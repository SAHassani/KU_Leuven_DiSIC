-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��V������6�8�!�%�+���Y����\��}��U���0�8�;�x�w�/����Ӷ��Y��N��<���c�`�_�x��)�M��Y����Q��^����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��Yۅ�V��-�����=�u�4�<�9�1�>�������G��X�����:�_�x��;�����Y����A��=C�;���:�4�u�;�#�(����Y����A��'�����!�:�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9K�g�����u��6�4�2�;�����Ƹ�VF��V�����u�0�<�4�8�s�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=d�����,���y� �/�L�������v#��D�����6�d�c�{�;�f�Wϫ�ӯ��vH��Z�����1�4�9�_�w�.�W���ݶ��u��C*��6���3�6�0�!�y�1�L�������VF��P(�����;�9�0�<�6�2�W���s���3��V�����&��6�0�2�)����
����G6��D��ʓ�4�!�0��8�����������=N��Xʼ�u��8�=�$���������@l�T�����u��8�=�$�����Y����T��S��F���x�u�g�{�e�}��������X(��t��%���0�<�&�o�>�)����C����F�=�[��u�6�;�!�9�}�3���6����]��T�����0�u�h�a�l�p�$��I���F��X��U���!�0�;�8�2�}�Ͻ�����Z��DN�����0�u�;�0�4�}��������r%��X�����x�1�6�8�#�2�W�������UF��=N��Xʾ�:�3�u�u��(��������R��X��U����8�4�&�~�r��������9F�N��U���u�u�� �3�-�E��Y����F�^�U���{�m�u�x�w�5�W�������@%��T-�����<� ��0�>�g�W��Y����Z��\-������-�0�<�6�4�������F������}�{�m�d�~�`�F��s�Ư�]��Y��8���4�6�,�9�$�g�������F�� UװU���u�=�&�!�'�}�ϫ��Ƹ���V�����,�u�3� �$�:��������G��^�����7�!�"�1�?�.�ϼ�s�����Z>�����!�_�u�,�2���������Z��E��]ʻ�!�'�9�'�9�8�K���Y����]��Y������4�0�<�$�l��������l�C��U���4� ��,�#�4�W������]��E�����0�k�|�:�w�4��������|��R �����d�1�"�!�w�t�}��� ����]��Y��4���!�<�u�'�6�u��������R��R�\ʺ�u�;�<�;�3�e��������l�C��U���;�1�m�'�e��W���������B��U���2�u�k�y�9�)��������Z�N��U���;�1�d�u�8�3���B���F��B�����&�;� �<�$�4�W��� Ӑ��Z��CN����&�:�9�u�2�<�ϫ�����V�N�U���;�<�2�!�>�}����Y����WF��F��ʷ�&�u�:�3�>�4��������G��B���ߊu�x��u������Y����T��V �����%�4�0�!�w�2�Ϫ��ƥ���SN�����!�_�u�x� �/�W���Y����VF��X����� �<�&�_�w�2����Ӎ��^6��T�����;�!�u�u�9�8����D����9F�N����� �6�<�;�w�8��������A����ʡ�0�'�2�!�$�?����ӥ��U ��E�����x�3�'�0�4�}����
����3��C@ךU���6�<�;��#�2��������R��t������&�4�6�m�4�����ƾ�G��,��8���!�_�u� �4�4�ϙ�����\��u��4���,�>�:�3��0��������Z��P��U��� �;���d��L����Ɯ�P��RN�����6�<�;�9�2�4����B���P��RN�����>��4�!�8�<�3���������=N�� ���<�;��!�8�;�5���8������R�����&�4�6�o�>�)����Y����A��e/��C���<�_�u�u�6�4����+����]'��V��U����c�!�o�w�2����Y���\��E��K��r�|�_�u�2�4�}���Y����p	��Q#��<���4�6�u�u�~�)��ԜY���a��E �����o�u��0�1�8����B�����^��6���3�0��&�6�>�W���PӒ��]l�N��'���'��'�,�m�}�4�������A��=N��U���0�u�u�u��)�������F��X��8���'�g�_�u�w�3�W���s���A��E �����;�'�4�n�w�8�ϙ�����U$��Z/����_�u� �6�>�3�0�������U ��V�����>�:�3��:�3�����ƥ�G��EG�����;���f��}����YӐ��Z��RN������'�,�o���Dف�Y���\��E��K���!�0�&�h�w�m�^��Yӄ��ZǻN��¾�:�3��8�9�)����D���G��=N��U���0� �;�'�6�}�Jϵ�����V��N/��E�ߊu�u�9�<����������G��RN��D���=�;�u�u�w�����8����\�\-�����8�'��!�l�}�Wϻ�
���F�e�����'�,�o�u��8��������GT��N�����<�n�u�u�%�)��������r��NUךU���u�0��!�8�;�5���8����l��SN�����0�7�1�u�<���������V��V��N�