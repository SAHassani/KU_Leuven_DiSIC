-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B%��Q#�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������4ǶN����g�u�0�0�5�/�E��s��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�}�|�e�l�W��� ����GF��C�����;�!� �0�#�}��������]l�/��U���=�&��&�%�8�}��7����]��~ �����;�&��!�%�<�W�������Z	��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�'�������g�������;�u�8�9�:�3�Ͽ�����d��_N�����u�0�%�u�>�)�����ƞ�^K��D�����u�8�8�'�y�6��������Z��X�����d�y�7�!�4�3����
����Z��EN��U���<�0�{�x�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���lǑ[�����<�0�n�u�"�8����W����_	��T1�C���9�n�u� �2�4��������P9��S@���ߠx�u�,�!�2�4�W�������V9��Qd�����,� ���l�(�ϋ�0����e��G�������_�x�$�3����
Ӓ��]��C�����;�<�,���8�:����ƥ�F��R �����u�>�:�3�>�)�W���Cӏ��Z��P��N���:�!�_�u�6�-����7���	F����*���<�n�u�&��8�3���Y�����D�����6�#�6�:�����������Y��E��u�&��0� �}�W���Cӏ��@��[���ߊu�&�4��3�}�W���Y����G��X	��*���!�'�d�1� �)�W���s�ƿ�p	��c�����o�:�!�&�3�1��������AN��X�����x�u�:�;�8�m�W������B%��Q#�����_�4�6�<�2�)����-�ƣ�#��X�����,�<�_�u�4�0����Ӵ�� T��dd��Uʲ�;�'�6�}�w�}�Wϗ�0����Q��A�����d�1�"�!�w�t�M���[����V��G�U���%�'�u�_�w�}�W���Y����@��B����u�u�u��w�}�ϭ�����T��=N��U���d�o�<�u�#��������F�v\��U���&�1� �:�>�f�W���Yӧ��	F����*���2�6�_�u�w�}�C���ƿ�W9��X	��N���u�u��o�>�}��������l�N��"���u�u�;�&�3�(����B���F��rN����!�
�9�2�4�f�Wϻ�Ӆ��C	��Y�U���#�:�>�&�0�)��ԜY�˺�\	��D���ߠu�&�2�4�w�.��������QF��D�����6�#�6�:�����������Y��E��u�&�2�4�w�.��������F��D�����6�#�6�:�����������Y��E���h�}�!�0�$�c�G���s����ZǑN�����&�_�u�:�w�}����Ƨ�\��^
��X���0�0�4�0�]�}�W�������a'��6�����u�x�=�:��}�9���!����V��LךU���x�=�:�
�w�>�ύ�����_��=N��U���=�:�
�u�w�.��������l�N����>�4�"�u�$�2����Y�����X��U��&��8�1�%�m�}���Y�˺�\	��VN��U���4��1�}�~�}�W������l��N��R���u�x�#�:�<�<����I���F�A�����4�u�e�_�w�}�Z�������\F��s��:���:�7��_�w�}�6��!µ��4��\��&���u�u�2�;�%�>����Q���F�'��!��u�w�e�e�g�m�^���Tӏ����h�����f�u�:�;�8�m�W��!����V��LךU���u�:�!�8�'�u�W���Y����F�
P�����4� ��8��t�W��Y����@��B���ߊu�u�u�u�g�}�J���
����W��G�U���u�x�<�u�$�9�������F�N��U���k�&��8�3�/�F��Y���K��YN�����9�2�6�u�w�}�Wϟ�Y���A��N��U���u�u�u�u�z�}��������\��=N��U���u�f�u�h�w�m�[���Y���F�N��Xʼ�u�&�1� �8�4�}���Y���rR�S�R��u�u�u�u�w�}�W���Tӏ����h�����u�u�u�u��}�W���
����U"��VF��Y���u�x�u�;�w�)�(�����ƹF�N��6���h�u�4�%�2�1�9��Y���K�^ ����� �:�<�_�w�}�W���<���F��t��"���u�u�u�u�w�p����
����_	��TdךU���u�0�0�4�2�����
��ƹ ��V��O���%�:�0�&��0�������F��P��U���<�u�<�<�0�8��������p
��OG�����u�u�u�&��)�8��������V�� ���8�n�u�u�2�9���YӃ����T��U���4��n�_�w�.��������[��D*������9�_�0�3��;��