-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��b�����&�&�{�=�]�p�6�������R��u�����<�=�&�7�#�3��������VF��X�����u�:�"�,�z�}��������A	��T�6����u�0�!�9�W�ZϚ����)��X��U��f�x�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���N��\�Fʖ�%�'�2�!��)����Y����A��Y��6���:�4�<�;�z�}��������4��R�����u�4�<�;�;���������/��R��ʜ�3�'�4�<�9�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǶN��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�x�_�x��/����Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���T���6��y�����<�&�&�u�>�1��������\��T�����u�0�1�1�1�3����
Ӓ��GF��RN�����x�_�x�%�8�4���� ӯ��vF��T�����u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W��s���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��X���u�=�u�,�2���������\��DN��U���0�u�:�8�#�5����7�ƿ�J
��P�����0�u�u�u�w�p�Z���������D��ʺ�u�=�u���.��������P��D��ʴ�1�&�6�u�w�$�ϼ����F�=C����;�8�u�&�;�6����Ӏ��_	��C�����!�;�u���-�����Ʈ�\
��Y1�����{�u�x�_�z��ϰ��ƻ�]A��T�����"�!�u�=�#�;����Y������,������6�:�w�>�}�W���Y���K��E�����4�2�:�u�?�4�ϸ�Ӓ��GF��V��U���:�u�u�u�w�}�W���Y���F�N��U���x�x�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W��T�Ƙ�VF��Y�����&�7�!�0�9�?����Ӈ����h�����'�u�:�!�8�8����Y����VF�N����r�r�<�u�8�}��������JF��S�����u�:�8�4�w�)����Yӵ��P��T��ǽ�2�u�u�u�z�W�Zϲ�����@F��E�����;�!�4�u�4�4�²��ƻ���^
��U���8�>�u�=�w�}�W���Y���K��C�����0�=�2�u�8�+�����ƹ�VF��RN�����0�u�4�0�w�)�(���������N��U���u�u�x�x�w�)�(���5����H�c�����#�x�:�u�2�.��������[��X��U���0�u�u�u�w�}�W���Y��ƴF��X1�����;�6�<�0�8��Wχ�Ӌ��[��E��ʡ�u�;�0�!�#�8��������VK��P��U���_�x�'�&�;�.����0ӕ��T�������=�u�6�<�2�1� Ͻ�����V��D��ʡ�0�<�!�;�w�}�Z�ԑTӏ��E�������!�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�C�X���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�z�p�W�������R��'��ʢ�<�!�;�w�2�4��������\��Q�����9�2�6�#�4�2�W������KǶN��ʹ�>�u�=�u�"�8�����ƾ�@�������;�3�'� �$�:���Y������V�����u�x�_�x�>�}����
������h�����0�!�'�<�w�2�W�������]F��D�����<�4�,�;�:�8�Y���T���1��X��ʢ�;�u�:�/�%�}����Ӓ����_�����4�u�3�9�1�q��������V��N��U���x�u�;�!�2�0����W�Ƙ�VF��XN�����:�&�w�0�8�����[����F��RN�����0�u�:�u�w�}�Z��Y����VF��V�����0�y�0�%�4�<��������A��^ �����4�9�u�0�>�)�������F�CחXʦ�8�u�;�&�3�?���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�x�]�p�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���l�������4� ��#�}�W���&����P9��T��]���1�"�!�u�~�}�W���Y���F�N��U���u�x�x�u�y�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���T���`��B�����h��'�&�f�t�Qϗ�����C��V��U�����$�0�#�{�8�������A��N��X�߇x�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�p�}��5����Z��Y�����!�u�0�%� �4�Ϭ�T����_��X�����&�u�=�6�w�(�W���Y���F�d�U���8�9�u�:�:�3�W���Ӓ��*��N�����:�u�;�!�2�-����ӄ��JH�N��U���u�u�u�x�z�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���9K�~N�����!�0��4�;�/����5����AF��Y�����8�2�!�'�6�2����Y����R
��SN�����x�_�x�4�3�����,����G��C��Yʡ�0�3�;�!�8�}����4����\
��S�����u�=�u�8�9�}�W��s���^��C��U���<�0�u�;���$�������C��V	��Uʁ�u�&�u�u�>�}�������Z�N��X���u� �!�7�w�<����[������SL��ʼ�u����0�4��������@��^ ��Y���u�u�u�u�w�}�Z�ԑT���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�1���� ӯ��v]ǻ��U����&�1�9�0�>�F��W����9F��D��0���;�8�'�6�$�9����s����X��>��;���<�<�<�&�$�}��ԜY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�U���u�&�3�9�6�/�Ϫ�	��ƹK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�!�%�w�2����/����AF�������u�4� �4�w�<���Y�ƣ���[��N���!�%�u�;�2�8�!����ƥ���V��U��� �4�u�4�0�}�I���ӏ��V��d�����u�4� �4��>����
Ӈ��R� �� ���u�4�2�u�i�}�ϰ�����l�C��U���f��,�!�>�}����Y�Ƣ�G��[N�����i�u�u�3�$�9��������G	��_�����:�e�n�u�#�-�W���Hŧ��l��DN�����}�;�!�'�;�/����E���\ ��C
�����
�0�!�'�f�}�������9l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�x�w�$�ϝ�����Z	��Q�����&�u�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s�����^�����u�:�#�'�>�3�W��Y����A��N�����:�u�:��8�8����Y�ƿ�W9��X	��\ʧ�!�'�u�:�;�<�L�ԜY����P��RN��ʶ�;�0�&�:�{�z�P��Y����9F��B �����!�
�:�9�6�����5���@F��D�� ���<�|�'�!�%�}������ƓF������=�2�u�:�!�/����Y����K������4�&�|�u�1�3����Y����\	��V �����}�u�u�!��2��������F��C��U���9�4��6�8�f�}���TӇ��Z��_��U���#�'�<�;�w�l�U��Yۀ��@�C��\���3�;�!�:�w�2�5�������P��v�����"�&�o�&�3�1��������AOǻN��U���u�u�u�u�w�}�W���Y���F�N�����;��:�0�9�8����s���F��C��U���=�6�;�0�$�2�[Ϫ����A��=N�� ���<�;�!�
�#���������\	��V �����'�u�!�
�;�:��ԶY���R��A�����:�#�'�<�9�}����Y���Aǻ�����;�!�
�!��:��������DN��N�����;�u�0� �9�.��������9l�C�����0�=�2�u�8�+��������A�������x�u�d�w�w�;�����Ƹ�l5��{�����!�'�7�o��2��������F��C��U���
�:�<�
�2�)��ԶY���R��A�����6�;�0�&�8�q�_����ƪ�_��C�W��_�u� �6�>�3��������Z��T��4���#��"�7�m���������\�N��U���u�u�u�u�w�}�W���Y���F�N��U��� �;�&�1�;�:��������9l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�x�w�4�ϸ�����]ǻC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u�z�}�����ƭ�@��[�����6�:�u�<�?�����Y����F��[N��ʡ�u�e�_�u�"�>����#����*��P��Oʻ�!�'�9�u�2�(�ϭ�����Z��R���ߠu�x�u�0�"�3�W�������T��A�����<�=��;�#�}����Y����@��C��D�ߊu� �6�<�9���������\��V�����'�!�'�u�#�����&����\��=N��Xʧ�!�'�&�6�>�4�ϱ�Y����T��X	�����_�u� �6�>�3�;���Q����	F��D�����'�!�'�u�6�(���s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�<�0��0�����ƪ�]��X ��U���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�W������]��_�����'�:�u�=�w�*�W�����ƹ ��T��ʙ�'�0�}�y�w�}��������V��YN�����'�_�u�x�w�<�W�������R��_�����!�u�4�9��/���Y���r
��DN��U���u� �%�'�2�}�ύ�����Z�� @�U���u�;�:�8�9�}��������W��V�����<�u�=�u�"�(����Tއ��R��V��ʙ�'�0�u�<�#�:��������AF��C��U���0�0��_�w�p�W�������G��D�����:�u�=�u� �}����
����F��^��&���9�'�4�7�m�4�����ƾ�G�������n�_�u�x��3��������AF��NN��U���9��4�9�%�}�?������D�������u�<�y�,�"�}�Z�������@��_�����1�1�;�8�w�
�%�������G��C��1����;�-�,�u�)�W������K��X�����&�"�!�u�?�}��������\��X�����!�&�u�0�>�8�W���Y���`2��d�����{�u�4�9�9�}�����ƥ���U��ʦ�8�9�'�_�w�p�6���
ӏ��]	��D�����1�7�u�,�'�4����N��ƹK�b �����!�!�0�4�>�.��������\��YN��ʳ�!�'�_�u�z�1�����ƥ�5��[��U���!�2�'�u�9�8����������R	��(�ߠu�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z���T�ƚ�P��/��Z���3�;�!�:�$�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǑN�U���&�u� �6�>�3�W�������[�x<�����#�'�u�<�w�;��������AF��D��U���u�3�;�!�8�}�������R��N�����2�6�#�6�8�t�����ƿ�W9��X	��N���3�;�!�:�w�/�����έ�TF��B �����|�'�!�'�w�)�(�������F��Y�����'�0�!�'��/�W�������]0��C��U��� �;�7�:�2�3�}���T�Ƙ�V��Q�����&�'�!�'�w�5�W͟�=�ƣ���E�����3�!�0�#�4�2�W���
����]l�Q�����u�;��6�8�}����Cӕ��l
��^�����'�u�0� �9�.��������9F��B ������1�0�!�%�u����Y����T��N�����u�!�
�9�0�>�}�������\��Y
�����u�4�2�o��2��������F��C��U���9�4�n�_�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F�=�����,��;�=�$�.�6�������@l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u�#�/����Y����[��T�����2�_�u�!�%�?���� ����R��U��Oʷ�:�0�;�_�w�)�����ƿ�]9��T�����u�!�<�2�]�}��������@��R ��*���:�<�2�o�$�/���YӇ��A��C�����0�%�o�7�8�8��ԜY����Z��RN�����'�6�
�;�5�8�Mϼ�����l�V�����0�&�;�8�/�<�W�������A]ǻ�����!�u�6�%�8�.�Mϭ�����9F��C�����u�,�
�:�;�>����Cӄ��_��d�����<� �0�9�4�����Cӕ��Z��=N�����7�!�u�,��.���������[��N�ߊu�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}���T�Ɗ�]��X �����&�!�<�2�5�)�X�������Z��YN�����:�_�u�x�w�1�W������� ��T�����0� �;�4�$�9��������G	��@��U���4�2�u�3�w�p�Wǉ�Hӂ��]��G����0��1�3�"�)�W���J�ƥ���^�����%�6�3�0�y�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǑN�U���8�9�&�_�w�p�W��Y����A��]����#�6�:�u�>�5����Y���J��Y
��Mʦ�!�u�x�u��>�E��Y����Z��[�D���d�|�n�u�z�W�W��7����VF��V�����4� �4�u�%�<�W���ӄ��V��X��U���%�'�;�=�$�.�W��� ��ƹK�Z��U���0�1� �9�w�<��������J	��T��U����!�{�u�2�8�Ͽ���������U���u�0�u�=�w�<�Ϭ�
����G�������4�0�!�0�%�<�����Ƹ�VF��C�����;�_�u�x�:�/�W�����ƹK�\8��F���h��!�<�$�����
���F��N�\��u�x�_�u�z�����Y�����������"�!�u�<�$�o�W��O�ƭ�WF�������x�>�0�c�w�`�$������J�N�U��y�c�|�_�w�p�WϿ�����G��[ךU���>�0�c�u�j�����
ۯ��Z��
P��Y��u�y�c�|�w�`�A���s���9F�N�����u�u�g�7�#�+����Y������]���ߊu�x�>�0�d�}�Jύ����� O��N����x��!�'�w�}�Eϼ�Ӑ��G	��@��U���u��7�<�w�<�����Ƹ�VF��[�����u�<�;�9�4�1����;��ƹK�V �����>�:��!�#�6����Ӓ����B��ʴ�&�2�4�u�6�1�Ϧ����K��a��G��u�0��!�<�2�5���Y����F��=��7���>�:��!�w����Y���F�<�� ���4�f�x�<�w�8������������ʼ�u�0�u�:�/�2�W���Y����K,��q��ʣ�6�:�u�&�w�p�W���������C�����u�!�'�<�0�<�W���Y����9F�N����u�h��!�>�u�5�������q	����&���<�9�}��2�}�=�������l�CךU����!�u�=�#�%��������R��RN��U���0�0�y�4�w�3�����ƣ���C
�����
�0�!�'�]�}�Z���T�ƀ�GA��D�����4�0�4�'�6�<��������V�&��ͦ�!�0�:�1� �$����ӏ��9F�d��X���'�6�&�u�:�2�[ϳ�����_�Z'�����;�_�u�x�5�:����T���^0��\��H���!�0�&�h�w�m�^�ԜY�����e�����!�1���0�}�>���������Yd��X���u�u��6�e�6���������UUךU���u�u�8�0�d�u�=�������@��X��ʾ�:��0�1�w�`����?����l�C��U���u�3�_�u�z�8�Ϯ�����l�CךU����1�=�'�p�}�����ƻ�J\ǻC�U���u��6�g�k�}����ۍ��Q$��N�����:�u�0��2�9����?����F��X�����_�u�x�u�w�}�W���Y�ƻ�V��R	�����0�}�,�0�{�0�������V
��F�����u�k�r�r�l�}�Z�ԜY����[�������;�u�'�u�;�2�����ƥ���C�����u�=�;�"�>�4�Ͽ�Ӕ��W��=N��Xʧ�2�&�0�&�w������Ƹ�VF��SN���ߊu�x�u�x�w�<���Yۉ��V��
P��E���_�u�x��#�u�5���Y���A��N�U���4�>�:��2�9����������R(�����u�x�u�u�w�}�W���Y���@��[�����6�:�}�:��.����Q����y	��^��&���|�n�u�x�w�/����)����~��PB�����n�u�x�_�w�p�6�������[��R����u�x�_�u�z�
��������+��R	�&���<�}��7�w�/�$�������X,��q�����l�|�_�u�1�3����Y����Z��~ �����o��!�'�;�8����Y����]��E��O���g�u�0� �9�.��������V��EUךU���6�<�;��#�4�_�������]��E�����u�u�u�u�w�}�W�������@��[����u�d�n�u�w�}�W���Y���F��T�����4�u�h�f�~�/����Y����_	��T1�����n�u�3�;�#�2�W���;����]��T�����4�n��o�9�)����C����F��C��U���
�:�<�
�2�)��ԜY����G��=��7����1�-�o�9�)����s���F�N��U���u��9�o�5�2����s���F�N��U���u��o�;�#�/���Y���A��E �����:�<�
�0�#�/�}�������\��R������1�-�o�9�)����s���F�N��U���u�u��9�m�(������ƹF�N��U���u�u�u�u�w�}��������U���� ���&�1�9�2�4�+����B����F��^��&���<�9�}�;�2�}�W�������9F�N��U���u�u�u�u�w�<�W�������T��A����u�u�u�u�w�}�W���Y����\��V�����h�f�|�'�#�/�W���&����P9��T��N���3�;�!�:�w�8�1���ۯ��V� �� ���n�u�u�u�w�}�W���Y���0��T�����4�n�u�u�w�}�W���Y���F��T�����4�u�h�f�~�/����Y����_	��T1�����n�_�;�u�6�6��������G��C��1���_��6�4�2�?��������G��C��1���<�_�u�x�w�5�W���ӕ��R��NN��U���u�:�#�'�2�}��������G��DN��U���"�<�0�:�2�}�Z���Ӓ�� ��T�����=�!�1�3�9�}��������\�/��U���u�!�0�u�"�>����s�����^ �����'�7�=�#�8�}�Ͻ���������ʳ�;�!�:�&�]�}�Z���T�ƅ���DN�����!�
�:�9�6�}��������	��TN��ʡ�0�7�&�u�"�>����W���F��RN�����u�:�#�'�2�.�����Ư�_
��_�����3�;�!�:�$�4��������l�C�����6�<�0�9� �>��������^��[�����!�!�0�'�$�1�ϱ�Y����Q��=N��Xʳ�;�!�:�&�]�}�Z���T�Ƙ�Z��G�����%�:�4�9�w�8����Y����R��Y��ʶ�1�y�7�!�>�}����Y���P	��R �����u�=�u�0�6�4�Ϸ��ƭ�@��[N�����u��u�=�w�4������ƹK�T�����'�u�'�u�8�/�������Q�������#�6�:�u�8�+����
Ӈ��9F�N�����u� �'�;�2�9����������C�����4�<�;�7�#�3�Ϫ����F��Y�����&�!�0�&�;�8�Y�ԜY����V ��RN��ʷ�&�u�:�#�%�4����T�ƙ�_����U����1�3�;�3�W�W��YӀ��P��YN��*���}�u�u�!�"�2�������	F��CG�����;�7�!�_�w�p�8�������A��
��ʻ�!�4�9�"�6�$��������G����U���u�4�0�"�2�W�W������]����U���0�4�#�9�2�}�?�������F�������&�;�u�:�%�>���YӀ��P��YN��*���9�4�u�&�m�.����������B�����0�;�<�_�w�8��ԜY�ƾ�G��F��*��}�|�r�r�l�}��������\
��YUװU���u�u�4�0�4�3����ӄ��V��YN��U���&�<�2�:�2�<����[����l�Q�����u�:��:�2�3�����������*���2�6�u�0�"�3��������@l�U�����u�'�!�'�w�	�(��Q���A�=N�����:��:�0�9�>������ƓF�/�����4�<�0�6�9�8������������ʶ�;�0�!�'�w�;�����Ƹ�l$��[��#���:�}�u�u�#�����&����\�E�����:�9�4��4�2�W���Y����R��U�����u�u�:�9�6�����Q����]��d�����;�u�u�3�%�4��������R�������u�u�'�4��t�M�������_����\��u�u�0�1�;�2�L���YӔ��F��E��N���0�1�!�
�8�1��������9l�C��U���<�4�<�0�4�3����ӓ��]��YN�����;�u�%�'�#�/�_Ͱ���ƹ ��T��ʡ�
�:�9�4��>��������\��T�����:�<�
�0�#�/�}���Y���F�N��U���u�u�u�u�w�}�W���Y����A��X�����6�:�u�&�w�}��������A��T�����4��6�:��z����P���Q��Yd��Uʳ�'�<�<�u�!�1����ӊ��Cl�N�����}�|�o�u�8���������E��@F�����_�u�u�;�w�2��ԜY�ƾ�G�����ߊu�;�u�:��2��������r��A���ߠu�x�u�=�w�<�Ͻ�����Z	��N�����:�u�:��3�2����Y�Ʈ�\
��YG�����;�&�1� �8�4�W���Yӄ��ZǻN��ʷ�!�0�_�u�w�}��������l�N���ߊu�u�u�0�"�3�P���s���V��^�Uʰ�1�!�
�!��:��ԶYӀ��P��YN��*����2�6�6�>�8����Y�Ʈ�\
��YG�����;�&�1� �8�4�W���Yӄ��ZǻN�����;�;�!�!��)�;���ۄ�9F��Y
�����1�:�<��#�+�;���s����F��^�����!��2�6�2�)�Ǽ�CӤ��_��a�����'�!�'�u�#�����&����\��Dd��Uʣ�'�4�9�u�!�1�Mϭ�����Z��R��·�'�;�0�n�w�?����Y����\�������r�4�2�u�8�-�W���YӔ��_N��T�����!��2�6�5�4�^�ԜY�Ʃ�WF��X�U���'�!�'�u�!�1�}����Ƹ�l5��{�����!�'�_�u�1�3����Y����G��P�����'�6�<�0�8�u�W�������]0��C�����u�u�u�u�w�}�W���Y���F�N��U���u�'�!�'�w�)�(�������P����Uʷ�2�;�u�u�%�)�����Ƹ�l5��{�����!�'�7�n�w�8�Ϫ�&����\��a�����!�#��"�]�}��������i��DF�����u�u�4� �6�t�����ƿ�W9��P�����:�u�&�u�w�+�����ƚ�P\��C
�����
�0�!�'�f�)�W������	[�X�����k�r�r�n�w�?����Y����V��YN���ߊu�;�u�0�8�f�}�������\��Y��9���!�u�u�4�"�<�^Ϭ�����@��[�����6�:�u�&�w�}��������e����*���<�
�0�!�%�l��������F��F�����u�k�r�r�l�}���������B��#���_�u�;�u�9�.�}���T�ƀ�TT��R�����=�u�0�9�9�}�Ͽ�����F��P�����u��4�%�2�<��������	l�CךU���0�!�!�u�"�}����T���T��E�����x�u�u�"�3�5�MϷ�����\�\ךU���u�|�_�u�z�}����Q���F�N����<�u�!�
�8�4�(�������Z��_�����:�e�n�u�z�}�W�������Z��Y�����9�2�}�<�#�t�FϺ�����O��N�U���u�:�!�o�8�)��������9F�N��\�ߊu�x�0�1�:�%�}�������\��X	�4���o�%�&�!�!�t�����Ƣ�G��[N�����u�4�<�7�2�����/�����B��N���u�#�'�4�;�}��������\��V����u�7�2�;�w�}�%�������\�UךU���=�3�0��0�g�W���T��ƓF�@��ʆ�<�!�1�'�w�}�W���	���F��_�����2�o�u�=�1�8�6���V����F�N������9�o�u�2�(����Y����9F���U���%�_�u�u�%�)��������e��=N�����:�g�_�u�1�3����Y����V����U���0�0�|�'�#�/�W�������Zǻ���ߊu�u�3�4�i�?����s���F��C��U��u�u�0�&�]�}�W���������N�����<�n�u�0�3�����B���U��C��U���9�0�}�y�w�}��������V��YN�����'�<�_�u�2�4�}���Y����Z�������u�u�'�!�%�}�L���YӃ��Vl�N�����'�u�n�u�w�8�Ϸ�B����]��Z����_�u�x��2�8����������B�����w��u�3�2�8�ϼ�Ӊ��G��A�����4�&�1�<�]�}��������A0��C��]���u�u�!�
�8�4�(������A��E �����9�2�6�<�]�}�W�������4��B�����u�!�
�9�0�>�}�������F�e�����9�o�u�e�l�}�Wϸ�ӏ��]F��PI�����9�:�_�u�w�}��������	[��R�����u�'�4�2�>�f�W�������\	��=N��U��� �;��!�%���ԜY����|��T��N�ߊu� �6�<�9��!�������A������1�u�0� �9�.��������Zǻ���ߊu�u�0� �9��!����ο�W9��P�����:�}�'�|�l�}����6����G	��=d�����!�:�u�'�2�)��������q	��R�����'�u�0� �9�?����ӏ��F��P��U���'�!�'�u�8�����۩��V��EF��*����2�6�0�#�/����P��ƹ��!�����'�_�u�x�w�5��������\��E�����=�u���w�;���� ӄ��	��C�����:�u�4�&�3�4�}�������\��Y
�����u�4�2�o�$�9��������G	���� ���&�1� �:�>�}����YӐ��Z��RN������9�o�&�3�(����B����V��=N��U��� �;�4�u�j�z�P�ԜY�ƪ�AF��^ �����4�2�u�:�'�}�W���+����]0��T��'���'��9�4�3�<�Ƿ�B��������ߊu�u�0� �9�����/����F��SN�����!�'�_�u�1�3����Y����V��EN�����u�;�<�;�3�}����ӕ��l��P���ߊu�0�<�_�w�}����ӧ��e��X�����:�<�
�0�#�/����P���V��v �����'�_�u�3�9�)��������G	����U���:�9�4��4�2�^Ϭ�����Q	��R���ߊu�0�<�_�w�}����Ӳ��q	��R��4���0�!�'���)�;�������\��E	��\�ߊu�;�u�;��>���s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߊu�x��;�#�2�ϸ�ӕ��G����ʴ�1�7�!�<�;�.� ����ƭ�E��XךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Z�������@F��D�����6�#�6�:�w�4�Ϫ�ӄ��@F��E�����<�2�!�u�9�4������ƹ ��T��ʆ�!�<�&��3�>���7����R
��T��Nʂ�o�;�!�'�;�g�W��Y����A��C
�����
�0�!�'�>�W�W�������_��V��Oʦ�1�9�2�6�!�>����T�ƨ�D��^����0�<�_�u�w�<���Yۉ��V��
P��E���_�u�u�:�w�}�ϗ�������P�����u�u�u��#�u�����Υ�F��I�N���u�0�1�9�8�f�W�������]F��C�Uʰ�1�3�;�!�8�}������ƓF�<�� ���u�u�!�
�8�4�(�������Z��U��<���-�u�0�u�8���������Z	��d�����;�0�u�u�6�(���Y���F�N��U���u�4�u�u�#�����Y���A��N��U���u�u�u�u�w�
�Mϰ�����\�\�����'�u�!�
�8�4�(�������@l�N�����9�u�4�4�m�.��������V��EF��Dʱ�"�!�u�|�]�}����s���K��Y�����!�4�&�4�2�2����YӇ��V��~ �����'�%�'�w���������Q��R�����u�w�&�#�%�)�W�����ƹF������<�u�'�;�;�)�(���Y����R��S�����'�u�k�r�p�f�W���=����z��OG��Hʃ�9�_�u�u�2�(�Ϛ���ƹ�������;��!�<�l�W�W��+����]����*���<�
�0�!�%�*�����Ʈ�GF��E�����<�2�!�u�9�8�W���W����F��^��&���<�}�;�0�w�}��������\��V�����h�f�|�'�#�/�W���&����P9��T��U���u�7�2�;�w�}�����Ɵ�G$��'�����1�-�u�6�`�P���Y����]ǻ��U���6�<�;��#�4�L�ԜY����V��Y��U���
�:�<�
�2�)�ϩ��Ʈ�GN��S��U���u�:��2�w�;�����Ɵ�G$��'�����u�4� �4�l�}�W���Y���F�N�����u�:�9�4�l�}�W���Y���F�N��U���4� �4�u�j�n�^Ϭ�����@��[�����6�:�u�&�w�?����Y����V��YN�����}�;�0�h��9��������\9��S"�����4�|�u�h� �f�Wϻ�Ӏ��P��YN�����n�_�u�x��)����ӕ��l
��^�����'�!�4�u�6�}��������V��Cd��X���=�u�<�u�8�4��������R����<���-�_�u� �4�4�ύ�����WN��S��Oʻ�!�'�9�_�w�}�W���Y���F�N���� �&�2�0�l�}�W���Y���F�N��U���u�4� �4�w�`�D�������]F��S1�����#�6�:�u�$�}�WϨ�����VF��C��U���
�:�<�
�2�)�ǉ�Hӂ��]��G��H���!�0�&�h�w�m�^�ԜY����]l�N����=�&�&�!�6�.������ƹF��D��ʜ�1�-�i��%�-����0������CN��U���&�!�4�u�u�.�����Ʃ�A	��=N��U���0�!�}�4�p�8����Rӯ��V�S�����u�u�0�:�#�����
Ӓ���������<�u�0�!�%�}��������A��d��U���&�;�=�&�$�)��������]l�N�����x�u�:�;�8�����Y����G��X	��*���!�'�'�&�-�u���.ޯ��V�d��Uʧ�!�'�u�4�6�W�W���Y����G��=��3���1�_�u�x�w�8����Y�ƿ�W9��P�����:�u�=�!�?�.�!�������]��VךU���!�0�7�!�'�.����Y����P��SN��U���0�{�u�3�9�)��������_��Y
��U���4� �4�n�w�}�W���Y���F�N�����u�!�
�:�>��������F�N��U���u�u�u��m�3������� T�E�����!�
�:�<��8�������Q��Yd��Uʧ�!�'�u�0��8�Ǘ����z��OB���� �&�2�0��<�^���Dͱ�9F��Y
�� ���<�;��!�>�1�L�ԜY����V��Y��U���
�:�<�
�2�)�Ϫ��Ƥ�@F��[N�����0�u�!�u�z�}�����Ƽ�@��X �����4�0�u�,��9��ԜY����G��=��3���1��1�-�m�3�������F�N��U���u�u�u��;�g��������F�N��U���u�u�u�u� �g�������F��N�����u�!�
�:�>�����ӏ��F��P��U���'�!�'�u�2�����0����X��S��U���h��
�;�>�3�ǈ��ƛ�z��OG�"���|�_�u�;�w�(����ӵ��u��SUװ����6�4�0�5�9�W���7����_��R���ߠ