-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��������!�:�o��3�5������|��^ ��U���?�6�o���p�A���s����R��_�1���8�0�u�e�e�p�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d�U¶�u�e�g��'�/����7����]��~ �����;�&��'�8�<����T�ƍ�_F��P��U���0�#�1�x�w�<����ӯ��G��R ��U���0�;�9��1�/�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�x�u� �'�.�M��s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߠ9�7�4�,�>�8�L�������V��D�����6�d�c�{�;�f�Wϫ�ӏ��VH��Z�����1�4�9�_��>����)������=N��Xʡ�<�u�4�4�#�-�W�������U	��G�����g�u�'�4�$�?����Ӆ��C	��Y��Uʆ�;�0�u�x�w���������@F��Q��ʷ�u�u�0�0�>�}�Ϫ�Ӓ��
��R�<͸�6�:�&�;�w�2����s�����
��ʷ�u�3�"�1�?�i�Y�������UF��X�����u�<�9�7�w�m�WǺ�	����]��Yd��X����!��1�?�}����	����I��X�����:�%�9�u�>�8�}��� ����C��C��U���4�'�,�}�9�8��������X�X�����:�<�
�0�#�/�C�������V�=d��X���=�&�1�!�w�$�Ϸ�Y���� �������u�=�u�4�'�8��������\��Dd�����u�:�;��4�)����������R	��U���2�u�k�u�1�(��������W	��C��\�ߠ0�1��2�&�W��������\��g��ʼ�_�0�1��0�,�}�