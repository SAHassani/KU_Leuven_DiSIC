-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����E��[�����,�6�:�;�2�s��ԑTӧ��[	��*��U���0�u�;�u�8�8�4�����ƴF��^	�����'�?�6�o���(��L���"��RT��Dʔ�2�&�u�e�e�p�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d�U¶�u�e�g��'�/����7����]��~ �����;�&��'�8�<����T�ƍ�_F��P��U���0�#�1�x�w�<����ӯ��G��R ��U���0�;�9��1�/�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�x�u� �'�.�Mϊ��Ư�^��R �����0�0�!�u�w�2����Y����
��DN�� ʦ�;�=�:�<�2�p�W���Y�����VN��U���4�!�'�6�8�6� ���Ӏ��B��T��ʴ�8�9�<�9�w�;����T���F�N�����&�:�<�<�6�}����W���F�N��U���u��0�6�8�6����Ӓ��@��^�����3�0� �;�.�/��������Cl�N��U���u�7�!�0�9�����Ӈ��)��E-��[���_�x�u�u�w�}�W���Y����A��XN�����=�u�#�'�;�>���� ����F��EN�����!�<�u�4�2�p�W���Y�����C�����;�0�;�9�$�<�����ƣ�G��D@�����4�u�:�1�5�)�������F�N��Uʴ�!�'�1�"�;�<��������c!��^��ʡ�u�0�%�!�>�}�����ƪ�\ǶN��U���u�u�:�2�>�:��������G��EN�����4�u�!�!�w�4����Y����_F��[N�����u�u�u�u�w�>����Y����@��[�!���u�0�!�'�w�.����Ӓ��R��SN�����8�u�=�;�z�}�W���Y����R��[��ʚ�0�6�>�6�:�}��������V��[��ʡ�4�u�4�u�6�8��ԑT���F�N�����u�!�'� �y�p�}��Y���F�X-�����$�4�&�e�6�}����������RN��U���0�9�u�;�w�3��������JF��C��U���u�u�0�0�.�����Ӆ��_�x �����0�4�!�'�8�2��������@l�N��U���u�>�#�'�;�>�1������J�� ��U���<�2�0�2�w�;�5���:����Z
��_�����x�u�u�u�w�}��������	��B �����&�7�6�u�8�m�WǍ�Ӓ��Z��S�����7�9�"�_�z�p�W���Y���	��B �����&�&�8�u�.�1�Ͽ�����a��CN��U���&�;�0�u�8�/����WӢ��Z��C��U���u�u�!�0�2�)��������P��R��6���!�4�<�u�$�;����Y����]��V��U���:�0�_�x�w�}�W���Y������YN�����u�&�&�;�2�}����������Y���߇x�x�u�u�w�}�Wϱ�����X#��R ��ʼ�u�'�0�!�2�>��������VF��RN�����u�1�0�:�w�<����W���F�N��U���&��>�1�2�8�Ͻ�ӄ��F�������;�7�0�&�0�<�W���Y����C��R��X���u�u�u�u�#�<�W����Ƹ���^��ʗ�&��>�&�0�<�Ϸ�Y����|��t�����<�u�<�=�]�p�W���Y���Q��E�����0�!��&��6�����Ʃ�T�CחX���u�u�u�u�?�}��������W��E�����&�'�!�&�#�8��������\�������:�>�;�u�6�)���Y���F���F�߇x�u�u�u�w�}�W���Y���F�N��*���
�u�u�u�w�}�(���&����F�N��U���
�
�
�x�w�}�W���YӤ��V%��N��Uʊ�)�u�u�u�w��(���&���F�N��*���
�
�u�u�w�}����&����Ol�N��U���u�u�u�u�w�}�W���Yӹ��F��hN��U���u�u�
�u�w��W���&���l9�N��U���
�_�x�u�w�}�W�������XF�N��*���)�
�u�)��}����YӚ��OF��h1��U���)�u�
�)�w�����&���9K�N��U���u�� �!�w�}�W��������N��U��u�u�e�u�w�l�W���K�ư�V�KN��Uʩ�u�u�)�x�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y�Ɠ�l9��h1��*���
�
�
�
���(���&����ll�N��U���u�:�:�;��1����&����l9��h1��*���
�)�x�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�(���Y���F�N��*���
�u�u�u�w�}�Wρ�&��ƴF�N�����9��2��/�}�(���&����l9��h��U���
�
�
�
���W���Y����l9��h1��	���u�)�x�u�w�}�9���CӉ��@��\+�����!�<�u�:�w�(�������G	��B��U���u�=�u�<�$�}��������Vl�N��U���u�u�:�:�9���������G�q�����%�0�<�u��8��������R��EN��Gʡ�0�3�'�!�z�}�W���Y���	��D�����0�0�!�"�;�}����Ӈ��V��t�����<�u�&�0�#�s�}��T���F�N����� �%�!�u�2�9�DϬ�
����V��DN��U���0�9�u�9�$�o�8���������[��X���u�u�u�u�6�)�Ϭ�
����V��R��U���&�;�u�'�'�/��ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C���7�4�,�<�2�f�Wϫ�ӏ��VH��S1�����d�c�{�9�l�}��������]��E�����4�9�_�<�%�/�W������F��@��[����%�4�9�]�}��������X��b�����&�&�{�9�l�W���� ө��A��T�����6�:�;�0�w�.�������F��A������6�:�u�w�g��������AF��]�Uʾ�:�;��-�6�2����Y����]F��E��U��w�e�|�_�8�)�}���+����F�N��U���u�u�o�<�w�2����B����R��[��U���u�u�u�u�w�}�ϭ�����Z��N�����u�u�u�u�w�}�W���Cӏ��Q	��R��O���'�0�_�u�!�/����Y���F�N��Oʼ�u�!�
�:�>�f�Wϱ�����F�N��U���u�u�u� �w�3����ۊ��
��D_��:���6�:�>�4�#�/�W������F��F�����h�r�r�n�w�2����/����F�N��U���u� �u�:�;�<�L�������p
��S	�����u�u�u�u�"�}��������V��x�����>�;��;��(����s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x��0�&�%�)����
ӕ��C
��=C�U��u�:�2�0�6��W����Ư�P
��^ �����4�0�9�u�8�<��ԑT���F��C��U���u�1�0�u�1�)�ϊ�����TF��d�U���|��9�,�#�8����Y����P��YN�����0�:�2�u�.�1�Ϫ�Y����V�������4�<�0�x�w�}�WϪ�Ӆ��]��N�����u�� �!�6�4�W���YӖ��@��u��6���1�0�0�!�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l��T�����'�u��u�1���������T5��T-�����u�&�u�&�0�<�W�������UF�T�����4�u�h�3�;�8�}���TӢ��V��Y�����<�0�:�u�?�}�1Ͻ����F�9�����u�:�4�:�3�1��������Z��C�����!�0�!�:�4�2�Ϻ�����F��X�����_�u�x�8�<�.�����Ƥ�A��XN������0�0�:�2�*�W���Ӈ��_��CN��ʓ�&�!�u�0�2�)�W��Y����W��^ �����:�2�<�2��s�Wϭ�����\2��P�����u�o�7�:�2�3�M�������9F��^	��ʺ�:�2�0��>�8�Mϼ�����\�Q���ߊu�x��0�#�}�W����ƞ�T��R��ʥ�%�9�;�u�2�<��������]��QN��ʰ�2�u�0�0�#�2�Y���T����VF��T��ʴ�u�0�&�u� �}����������V��ʺ�!�:�u�:�9�.��������Z��_�����_�u�x�'�0�.����
����^��d�����!�;�u�>�2�<�4�������\��Y�����h��'�0�w�o��������X ��C��N���&�2�4�u�w�2��������c��T�����4��6�:����������Z��N�U���;�:�e�_�w�}�W���Y���F�N��U���u�o�u�:�?�/�J�������l�C��0����!�6��'�u�^ϩ��Ƽ�_��X �����0�4�!�'�6�/����Y����	��u��6���_�u�x�:�6�8��������GF��X��U���&�u��0�4�2�������T��N��ʹ�!�'�u�=�%�;�������F��R
��ʱ�<�0�<�u�%�0��������P��G��:���6�:�>�4�#�/�Z��WӲ���������:�_�u�x�>�}�����Ƥ�]�������=�'�u��2�>����������[��U���;�f�_�u�8�.����Y����V%��r
��;����1�-�o�>�)����Y���F�N��U���u�u�u�u�w�}�W���Y���X)��E�����6�:�u�u�~�0�ϵ�����\��V���ߊu�x�:�:�9�}�Ϭ�
����V��Y�����u�,�9�u�1�8�W���
����v��y��U���&�&�_�u�8�.����Y����G��t�����0�u�u�o�>�)����Y���F�N��U���u�u�u�u�w�}�W���Y���X)��E�����6�:�u�u�~�0�ϵ�����\��V���ߠu�x�u�'�6�8����ӕ��]����U���%�!�u�0� �1�W���ӏ��Z��C��U��� �0�_�u�>�3����Y����]��[N��U���o� �&�2�2�u�4���Ԕ��T�S�����'�u�k�r�p�f�Wϭ�����F��t�����<��9�u�w�2����Y����R
��dךU����0�!�u�.�>�%���ӵ��]��d�����4�u�u�7�9�?����Y���F��U�����o�u�4�&�l�}���������V��U���u�u�u�o�5�2����C�ƪ�_��=d��X���=�u�#�'�;�>���� ����F��EN��ʷ�u�&�1�:�w�<�Ͻ�����]��V�����4�0�!�8�]�}�Zϭ���������ʖ�:�>�4�1��.�Ϸ�	����2��DN�����&�!�0�6�:�4�Ϫ�����RǻC����0�4�9�!�2���������T5��T-�����u�;�:�4�$�3��������V��V �����!�_�u�x�4�3��������F��C��ʓ�&�:�u�0�.�9����ӵ��P��X �������u�:�6�2����T�Ƹ�Z��RN��ʴ�>�0�u�!�%�?���-����D����ʦ�'�u�#�'�w�4�Ϫ����F��R�����;��;��"�)�Ϸ�Y����R��V��U���0�u�� �#�>�W�������V�N����� �0�>�0�w�}�������R��^��ʾ�0�u�3�:�8�3�;���Y����R
��DN�����n�_�u�x��0�W���	����G��D��6���!�!�u�'�!�}����	����Z��[�1���<�2�!�:�:�3�W�������F������9�6�;�u�9�}�����ơ�A��^�����{�u�x�u�?�}����������E�����9�:�u�4�?�4�����ƣ�)��E�����2�,�6�:�9�8�W���Y���P��D��U���<� �u�4�w�(�W���Y����]�N����� �0�8�-�1�3���
����T]ǻ�����!�u�4�
�6�2�ϱ�Y����]��[N����4�u�&�>�8�3�:�������l��R	�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}���T���p��C��U���2�0��{�w�5�Ϸ�Y������D��U���'�u�4�0�;�}�����ƥ���=N��X���u�#�'�9�w�2����Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߊu�:�2�0�1�W�W�������R4��R�7����>�u�&�w�?����Y����UF��R��U���;�u�u�u�5�3������� ��D�U���u�7�;�7�2�}�W������l�N�����2�0�3�u�j�;����s���V
��QN�����
�1�0��$�������ƹF������'�u�=�;�w�}�W�������_��DN�U���0�_�u�u�w�3�W���s���F��Y�����u�h�7�;�5�8���Y���K�`�����u�4�!�7�8�:�����Ư�R�������!�9�u� �w�;�����Ƹ���^
ךU���u�x�8�!�$�<���� Ӗ��Q
��D@ךU���u�3�7�;�5�8����s���F�U:�����3�i�u�:�w�	����?��ƹF���U���_�u�u�;�w�;�}����Ƽ�\��DN������n�_�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F�\��1���6�u�=�u�3�8�W�������\��^ ��3���u�x�u�|��1�Ϫ�Ӄ��VF��C�����%�9�0�0�8�:�W�������\F��X�����0�;�!�4�>�8�W��Y����[��X�����4�&�'�u��(�����ƭ�WF��B��U���&��>�1�2�8��ԜY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���� �!�'�]�}����
�έ�V��N�����>�u�&�u�5�:����Yӏ��R4��R�����u�u�u�:�8�:����Y���Z�Q���ߊu�u�u��0�1�1���	���[��V��N���u�u�:�1�2�8��������v��s�����%�r�<�=�3�*����P���	��R��H���4�&�|�_�w�}�W���
����v��y��U��3�9�0�_�w�}�W�������_F�N��H���!�0�&�h�w�m�^�ԜY���\%��Y�����6�u�h�3�;�8�}���YӃ��Z ��^�����2�}�#�'�;�t����s���F�:��ʶ�:�>�1�8�>�}��������[	��SN��U���1�0�u�'�'�/�ϼ�Y����k��YךU���u�x�!�:�$�}����
�Ƹ�V��E�����0�u�9�6�w�2����W���F��c�����u�u�u�h�5�2�������F�X:�����3�<�0�i�w�	����?��ƓF�N�U���&�1�u�=�$�-����
�ƣ�W��R�����0�e�u�h�8�2����Ӟ��	��P	��3���%�_�u�u�w�p�'���������R
��U���0�!�1�!�%�(�Ϫ�Ӊ��T��C��%���u��6�4�9�W�W���Y����V"��R�����:�1�0�0�2�)��������W	��C��\���h�:�1�0�2�8����ۉ��T��C��%���r�<�=�x�f�9� ���Y����9F�N��Xʖ�0�!�u�=�w���������}��N��U���9�7�u�'�2�2�����ƣ�VF��T��U���u�,�9�_�w�}�W������VF��RN�����4�0�9�u�>�4�ϻ���ƹF������>�1�0�0�#�a�W�������V��^�����0�9��2��%�>�����ƓF�N�U���4�0�!�0�4�(����Y����R��^����4�!�'�4�%�.��������UF��D�����u�u�<�u��:�3�������VN��R����� �!�;�0�~�)��ԜY���F��X��9���u�u�u�h��)����D���O��N��U���:�:�;��;�9����DӒ��V]ǑN��U���u�� ����6���)�ƣ�\��{�����:�u�!�'�w�0��������R ��EN�����_�u�u�u�z�9��������V��D��0����!�6��'�}����:����e��S"��U���u�4�&�u�?�1�}���Y�����P	��3���&�1�&�7�2�f����UӒ����Y�����&�'�&�!�>�}����s���F��D�����;��9�1�4�}����Y���F��t�����u�h�:�:�9�����H���F�R ����u�u�0�1�>�f�Wϻ�Ӗ��P��-�����n�_�u�x��)����Ӄ��VF��������{�u�:�3�8��������V�S�����2�0�3�-�%�2��������C�=d��X���&�<�;�!�2�2����
����p	��C8�����h�:�:�;��1����B����p	��CN��U���h�:�:�;��1�}���Y����9