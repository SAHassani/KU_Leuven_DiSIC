-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����9�6��%��s��ԑTӧ��[	��$��ʔ�8�'�4�_�z������Ɯ�\��CT��-���`�a��x�w�<����HӬ��JF��_חX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�������W��X�����u�4�<�;�;���������%��G�����_�x��9��:��������VǶN�����4�u�;�!�"�8��������R
��Y�����:�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s��ƴF��E�����=�&�3�9�w�4��������_��DN�����=�u�!�
�8�4�W����Ƹ�R��_חX���u�u�u�u����������(��RN�����0�u�:�!�2�3�­�����Z��X��U���!�0�x�u�w�}�W���?����w��E������%�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l��U��ʼ�0�y�"�'�l�}��������@��[����c�{�9�n�w�(�Ϸ��Ȣ�^��T1��Ĵ�9�_�u�&�w�2��������Z
��^�����9�n�u� �2�*����������d�� ���"�'�{�>��<��������Z��X����_�;�<�,��<����)����_	��c��9���&�u�2�;�%�>�}���Y����F��Z������6�0�o�>�}�����ƾ�]��N��U���h�a�_�u�w���������P��N��U��<�u�;�0�2�}����Y�Ƹ�U�
N����u��8�'�4�1����Y���F��^ �����0�u�4�2�w�}���C����l�G��]���u��8�9��6�MϷ�Y����_	��TUךU���#�'�9�u�w�3��������l�N�����0�0�u�u�9�.��������F�D+�� ���!��u�u�9�.��������9F������;�'�8�;�w�}�ϭ�����Z��R����u�:�;�:�g�f�W��H�ƥ�G��EN���ߊu�u��9��>��������VF��^ �����:�<�
�0�#�/�@Ϻ�����O��C��M��u�u�&�&��)����Y�ƥ���h����_�u�u��6�)����/����\��YN�����2�6�#�6�8�u�W������]ǻN��&���!�=�&�e�m�4�W���&����P9��T��]��1�"�!�u�~�}�Z�J����F�D=�����4�0�u�u�9�.��������V��EF�U���;�:�e�n�w�p�E���K�����V�����g�o�<�u�#�����&����\�N�����u�|�u�x��n�F�ԜY�ƿ�G��g�����u�;�&�1�;�:��������T��X����n�u�x�g�y�o�W���
����G6��D�Oʼ�u�!�
�:�>���������W	��C��\���x� �f�d�]�}�W�������R��T��ʦ�1�9�2�6�!�>����Kӂ��]��G�U���g�{�g�u�w�.����)����F��^ �����:�<�
�0�#�/�E�������V�N� ��d�_�u�u��<����
�����D�����6�#�6�:��o��������F�;�[��_�u�u��6�����
����Z��C
�����
�0�!�'�o�9� ���Y����K��@�U���&�0�1�1�%�.�F���ƿ�W9��P�����:�}�u�:�9�2�G��T�ƙ�_ǻN��'����1�0�&�w�}�ϭ�����Z��R����1�"�!�u�~�}�Zϋ�W���F��R�����&�f�o�<�w�)�(�������P��V�����:�e�n�x�w�d�N���Yӕ��R��S�����u�;�&�1�;�:��������F��@ ��U���u�x� �{�]�}�W�������A��N����!�
�:�<��8����Aӂ��]��G�X���l�l�u�u�$�8��������\��YN�����2�6�#�6�8�u�W������]�N��[�ߊu�u��4��9����Y�ƥ���h�����0�!�'�m�3�*����P���3��dךU����!���;�9�MϷ�Y����_	��T1�����}�u�:�;�8�m�L���Yӕ��G��~^��U���&�1�9�2�4�+����Q����\��XN�N���u�d�{�_�w�}�3���0����	F����*���<�
�0�!�%�l�W������]�N��M��u�u�&�4�6�3�E���ƿ�W9��P�����:�}�b�1� �)�W���Y����^�=N��U���!���u�w�3��������l��C��D���:�;�:�e�l�p�W��W���F��V����o�<�u�!��2��������W��S�����|�u�x��o�l�W���
����z��T��ʦ�1�9�2�6�!�>����Nӂ��]��G�X���d�{�_�u�w�����(����Z��C
�����
�0�!�'�f�}�������K�d_�D���u�&�4�4�9�n�MϷ�Y����_	��T1�����}�b�1�"�#�}�^���Tӵ��WǑN����� ��!�4�>�}�W���Y����_	��T1�����}�u�:�;�8�m�L���Yӕ��P��B��U��� �u�!�
�8�4�(������F��@ ��U���u�x�u�a�y�W�W���8����|��N����&�1�9�2�4�+����Q����\��XN�N���x��`�e�w�}��������zW���U���
�:�<�
�2�)���Y����G	�U��X���a�{�_�u�w���������	F��CN�����2�6�#�6�8�u�CϺ�����O��C�&���e�u�u�&�4�(�8���K����F��C
�����
�0�!�'�c�}�������F�=�[�ߊu�u��6�:�(�&���Y����@��[�����6�:�}�a�3�*����P���F��@�U���&�6� ��#�n�Mϱ�ӕ��l
��^�����'�a�u�:�9�2�G��Y����S�=N��U���6�8� ��w�}��������T��A�����a�1�"�!�w�t�W��Y����l�N������!�a�o�8�)��������l��C��A���:�;�:�e�l�}�Zύ�L��ƹF��v������u�u� �w�)�(�������P��Z����!�u�|�u�z�}�C���s���@'��B�����o�:�!�&�3�1��������AN��
�����e�n�u�x��h�G���Yӕ��P��B��U��� �u�!�
�8�4�(������F��@ ��U���u�x�u�a�y�W�W���8����|��N����&�1�9�2�4�+����Q����\��XN�N���x��`�e�w�}��������bP���U���
�:�<�
�2�)���Y����G	�U��X���a�{�_�u�w���������	F��CN�����2�6�#�6�8�u�CϺ�����O��C�&���e�u�u�&�4�(�8���N����F��C
�����
�0�!�'�c�}�������F�N��@��0�1��4�#�8�'���;����g	��{8����=�!�6� �2��;ϱ�Y����G"��g��7���>�:���>�W�W��Y����G��YN�����!�u�4�>�$�<����Y����R��NN�����&�u�x�u�2�8����ӄ��G��Z�����;�8�0�u�1��4ϭ�	����VǻC����=�u���]�}����ӕ��G��E�����u�<�;�1�o�/����Q�ƨ�D��^����<�;�9�&�6�<����0���5��Y��M���4�
�}�u�8�3���B����Z��[N������4�0�'�6�}�W���
����l�
�����e�n�u�&�0�<�W�������A��v���� �&�2�0�n�/�(���Y����G	�UךU���;�9�&�6�"���������"��V!��4���!�b�1�"�#�}�^�ԜY����R
��v������<�;�1�w�<����8����Q��X����n�u�&�2�6�}�6�������R
��u��Oʗ�:�0�;�0�#�/�@Ϻ�����O�
N�����&�h�u�4�$�t�}���T���E��\1�����'�_�u�x�z�+����
����Wl��R	�����x�u�4�>�#�8�3���0�Ɵ�eF��G��U���:�4�u�'�6�s�8���Y����U��Cd��X����%�!�4�'�8�'��� ����V
��R ��U���!�0�4�'�.�*����Ӆ��]��R
ךU���1�"�&�'�6�}�Ͽ�����]��R������{�u�&�6�<����0���F��^	��¦�4�4�;�f�{�}�W���Y���F�N��U���;�1�&�4�6�3�E��Y���F�N��U���u�u�<�;�3�.�������9F�N��U���u�u�u�u�w�4����
����z��G�����!��'�.�3�W��Q����V��s��<���|�_�u�u�w�}�W���Y���F��P ��]���!���|�]�}�W���Y���F�N�����0�}��!���^�ԜY���F�N��U���u�&�2�0������(���9l�D=�����4�0�'�4�w�a�Wǫ�
����WN��C��%���0�|�_�u�w�}�W���Y���F�N�� ���2�0�}��6�)����O��ƹF�N��U���u�u�u�u�w�}��������`��C>�����y�u�u�u�w�}�W���Y���F������1�&�!�'��<����s���F�N��U���u�u�u�u�"�.����Q����A��V��\�ߊu�u�u�u�w�}�W���Y���F��D������4�!�=�$�o�[���Y���F�N��U���u�u�u�;�>�3�ǭ�����[��G�U���u�u�u�u�w�}�W���Y����]��Y�����'��4�0�~�f�}���+����W��D�����i�u� �&�0�8�_�������A�� G�U���u�u�u�u�w�}�W���Y����]��Y�����1�1�'�&�a�q�W���Y���F�N��U���u�u�;�<�9�9��������V��BךU���u�u�u�u�w�}�W���Y�ƹ�@��R
��'����1�0�&�~�W�W���Y���F�N��U���u� �&�2�2�u�%���8����@��d��U���u�u�u�u�w�}�W���Yӓ��Z��SF�����1�'�&�g�{�}�W���Y���F�N��U���u�;�<�;�3�.��������@W�=N��U���u�u�u�u�w�}�W���Y����T�������1�0�&�|�l�W�W�������VF��V�����:��:�>�8�W�W�������RF��D�����u�u�u�u�w�}����������R�����_�u�x�=�8��W���6����G ��N��U���u�:�7�:�2�3��������u ��=N��X���:�
�u��6�8��������F������1�&�=�&��>�������K��X��ʦ�4�6�,�9�$�4�����ƹ�@��R
��6����6�0��9�.����Y����[	��h�� ���9��0�3�w�}�W�������\
��YF�����!�:�3�|�w�p��������`��C>�����9�1�u�u�#���������G	��D=�����4�0�4�<����������X�_�����:�e�|�u�z�+����ӕ��R��_��U���u�u�u�&�#�/�'�������JN��B�����:�>�u�u�w�2����I���K��X��ʦ�0�1�1�'�$�}�W���Y�ƿ�V��S
�����'�,�>� ��2�5������F��@ ��U���u�x�#�:�<�<��������_��N��U���!�
�:�9�6�����Q����R/��V��]���%�!�4�%�2��������F��@ ��U���_�u�x�=�8��W�������F�N��U���u��!��%�$����0����`��[�����6�0�x�d�3�*����P�����X��U���!���u�w�}�W���Yӕ��G��E������%�!�4�'�8�'��� ����F��S�����|�u�x�#�8�6�ϭ�����F��[��U���u�&�6� ��)����;����X(��g��7���>�u�u�u�8�3���s���E��\1����� ��!�u�w�}�W���Y����F��C'�����}��8�'�4�1����T����\��XN����x�=�:�
�w��������F�N��U���6�8� ��>�3�ǵ�����P$��T��X��1�"�!�u�~�}�1�������A	��[��!���o�0�!�!�w�2��������P6��T,�����%�}��|�w�}��������R�=N��U����8�'�6�;�>����Y���X��y�����9�6�&�u�w�}�W���Tӏ����R	��U���2�u�u�:�o�g�W�ԜY���X/��B�����&�0��6�2�`�W���	����^��D>��6���0�u�x�u�9�}�����ƾ�]��N��U���h�d�u�u�w�6��������R��EN��U���k�>�#�'�;�>�1������F�C����<�!�2�'�%�3�������	[�=N��U���!�8�%�}�w�}�Wύ�����_�N��U���u�k��8�;�����Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U�ߊu�u�u�#�%�1�W���Y���F�
P�����9�y�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���l�N�����'�0�0�u�w�}�W���D�Ƹ�l��[��]���0��&�!�{�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y����v��C��3���u�u�u�u�i�)�(�������@#��B�����|�u�u�u�w�}�W���Y���F�N��U���u�u�_�u�w�}�"�������U �N��U��u�:�7�:�2�3����8����V ��N��U���u�u�u�u�w�}�W���Y���F�N��U���u�&�=�&��>�������[�B �����}��4�0�9�/����P���F�N��U���u�u�u�u�w�}�W���Y��ƹF������6�0��;�$�3�W�������]��D-�����9�&�<� ��8�[���Y���F�N��U���u�u�u�u�w�W�W���Y����A��V�����u�u�h�u�8���������\��d�����&��9�1�<�(�'���;����@F�N�����u�|�y�u�w�}��������@�N��U���k�&�!�'��<�����Χ�F��X�����u�u�u�:�9�2�G��Y���F�N�����u�u��4��9����Y���F������1�0�&�'�6�u�9�������\��C��U���;�:�e�y�w�}�W���Y���F�N�����;�4�<�u�w�}�W��Y����\	��V �����}��!���1�ǵ�����R��R�����9�u�u�u�8�3���P���F�D*�����u�u�u�u�w�}�J���=����A��~ ����� ��8�9�$�8�4��������Y��E���u�u�u�u�w�}�W���
����z��N��U���u�u�k�&�6�<����0����z��C=������'�,�9�w�}�W������J�N��U���_�u�u�u��>����/����F�N��U���6�8� ��;�9��������A	��[�����d�1�"�!�w�t�W���Y���F�N��Uʦ�6� ��!�w�}�W���Y���@'��B�����2�0�}��:�/�������W��X����y�u�u�u�w�}�W���Y�����T�� ���u�u�u�u�w�c��������b5��Y������:��:�<�}�W�������V�N��U���u�u�u�_�w�p�6����ƃ�G��Dd����� ��!�4�>�}�JϪ�&����\��A������6�8� ��1������ƹ��T�� ���u�i�u�!��2����������T�� ���<�;�1�e�~�W�W�������G/��R�����9�2�6�#�4�2�_�������G/��P ��]���n�u�&�6�"����Y����G��X	��*���!�'�&�6�"���������O�=N��4���8� ��u�k�}��������E��X��4���8� ��<�9�9�D���s�ƿ�P��x��A���h�&�1�9�0�>�����ο�P��x��&���0�}�|�n�w�.����6����F���*���<�
�0�!�%�.����6����Z��SF�\�ߊu��6�8�"��W��Y����_	��T1�����}��6�8�"��������l�D/�� ���!�b�u�h�$�9��������G	��D/�� ���!��2�0��t�L���
����^)��f^��I���!�
�:�<��8����
����^)��f=�����e�|�_�u��>����(���F��S1�����#�6�:�}��>����(����V�G�Uʦ�6� ��!�e�}�Jϭ�����Z��R��¦�6� ��!��:����P��ƹ��T�� ���u�i�u�!��2����������T�� ���<�;�1�f�~�W�W�������G7��R�����9�2�6�#�4�2�_�������G7��P ��]���n�u�&�6�"����Y����G��X	��*���!�'�&�6�"���������O�=N��4���8� ��u�k�}��������E��X��4���8� ��<�9�9�A���s�ƿ�P��x��B���h�&�1�9�0�>�����ο�P��x��&���0�}�|�n�2�9�%���s