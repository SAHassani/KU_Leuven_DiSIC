-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s����c�:�9�#�3�p�W�������y	��-�����_�x��<�>�<�W�������6��R1�A܇�x�u�4�0�w�n�:���K����KǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��t�E��Y����A��CN�����4�u�;�!�"�8��������R��Yd�U���u�<�=�&��.����s����R��Y��<���'�8�;�&��)����Y����A��^��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��)����@��:��ʳ�9�u�&�&�4�<����*����#��C�����0�4�&�9�4�<��������]��R�����u�u�u�u�w�;����Y���^��N��ʳ�'�4�7�:�2�3������ƴl�N��U���u�u�=�u�"�-�ϭ�Y������NN��U���u�;� �u��9����ӄ��K�N��U���u��%�9�9���������[��E��U���9�&�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l��U��ʼ�0�y�"�'�l�}��������@��[����c�{�9�n�w�(�Ϸ��Ȣ�^��T1��Ĵ�9�_�u�&�w�2��������G��V�����!�'�4�9�]�}��������X��b�����&�&�{�9�l�}��������c��D����_�<�'�'�w��$���s�ƹ�VF��~=��[���8�:�0�!�y�1�L������� ��T�����g�c�:�9�>�W�W������F��Z��6���o�<�u�!��2���s���K��^�����1�9�,�<�w�$����s���@6��R�����4��;�&�?�8�W���ӓ��Z��SF����!�u�|�u�z��Y�ԶY���F��P ��U���7�u�0�4�2�W�W���=����]F��X���ߠu�u�x�u�>�3�Ϻ�����9F���Oʺ�!�7�:�0�9�f�Wϻ�Ӡ��P��T=��G���:�9�_�4�4�4�����ƞ�F��(�����6�'�g�c�8�1��ԶYӅ��C	��Y��'���g�_�u�u�8�)�_���Y����_������9�2�6�o�w�m�L���Y����\��YN�����2�6�o�u�g�f�W���YӅ��	F����*���<�u�h�r�p�W�W���Y����Z��C
�����
�0�!�'�c�9� ���Y����F�N��Oʺ�!�&�1�9�0�>�}���Y�ƽ�F��X�����9�2�6�n�w�8�Ͻ�����]��=dךU����u�0�1�6�+�����ƨ�_��Q��U���:�g�c�6�4�8�Yω�Y������[�����!� �<�2���E��Y���v��=��6���u�&�1�<�.�>����Ӓ��G��Y��U���y�0�6�u�;�0����Ӓ����^ �����x�u�0�4�2�}�EϽ�����^	����ʡ�0�%�0�<�"�}������ƹ��D��ʾ� ���9�e�g�������F��A�N���&�2�4�u��1����:����\��C
�����
�0�!�'�<�(�8�������\��XN�U��}�!�0�&�j�}�G���s�ƿ�T�������,�o�&�1�;�:��������X(��x����d�1�"�!�w�t�M�������@F�I�\�ߊu�<�;�9�$�/�&���)����	F��S1�����#�6�:�}��0����J����W	��C��\��u�:�=�'�w�c�P���B����Z��[N����� �3�1�9�w�}�������� ��D����x��9�!�2��;�������������0�{�u�&�0�<�W�������r��R��9���o�&�1�9�0�>��������W	��C��\�ߊu�<�;�9�$�/�:��������R	��U���2�u�u�:�9�2�G�ԶY���~����ʡ�<�u�<�;�;�4�W���Y����V��^�������u�0�8�8���YӇ��A��C�����o�&�'�;�l�}����������GN��U���!��3���$�Mϭ�����Z�C��W�ߊu�!�'�7�#�}�����ƿ�A
��E�����u�<�;�9�>�}����[��ƹK��_��*���&�4�!�u�z�+����
����Wl��P�����x��0�!�w�5�W���Ӌ��\��d<�����u�1�'�&�]�}�$�������W��D=��U��&�1�9�2�4�+����Q����V
��R*�����;�&�=�0����������V��{8�����|�n�u�&�%�����Y����\9��C��¦�<�0�<�0�2�<�:���
����VN��S�����|�n�_�u�z�����Ӓ����B��ʡ�0�3�'�!�������Ư�R��:��U���&�4�0�1�>�$��������@��=N��Xʤ�d�u�=�6�w�.�ϭ�����	��G�����=�u��u�?�)��������R�������4�0�u�:�#�}����T�Ƹ�VF��O��'���{�u�&�'��4��������Z�C�����2�6�&�|�]�}�0�������V��[]����:�u�u�;�<�(�8��������Y��Eʲ�;�'�!�_�w�}�Z����Ɵ�%��rN��'���g��u�u�z�+����Ӆ��5��G���ߊu�u�x�=�8��W���Y����w��N-�����|�u�u�x�!�2�������AǻN��X���:�
�u�u�w���������V��{8ךU���x�=�:�
�w�}�W��������N��Xǣ�:�>�4�$�f�.��������R��^E����u���g��}�%���K���F�G��U���u�_�u�u�w�}����Gӵ��C
��[�U���u�u�u�u�z�4�Wϭ�����Z�
N��R���u�u�u�1�w�`�W�������J%��^ ��\���u�x�u�;�w�)�(�������A��=N��U���u�0�u�k�p�z�W���Y���F�N��U���<�u�&�1�;�:���Y���F�N�����h�u��9�2�9����
����F�C�����!�
�:�<��8����Mӂ��]��GךU���u�u�u�u�i�.�����Υ�F�N��U���x�:�!�&�3�1����Y���F��_��Kʦ�'��<�,�?�4�_���P���F��CN�����2�6�u�0�3�:�����Ƌ�]%��T�����f�n�_�u�%�>��������p
��=N�����_�u�u�3�%�.��������R��R-��\ʡ�0�_�u�u�w�p�>����ƭ�u ��^	��U���!�0�#�'�6�1�W����ƣ�G��DN��U���u��&�u�1�)�����ƭ�JF��P��U���u�x�u�3�2�}����+����[��Z�����!�8�;�u�$�+��������F
��=N��U����9��,�>�8�K���*����A��=N��U���x��9�6�w�5�W���	����A	��C��&���!�4�u�4�w�5�W����ƨ�_��U��ʺ�u�!�u�:�>�4�Ϸ�s���F���U���<�{�u�u�w�.��������w
��S�����:�0�;�&�%�����	�ο�A
��O=��\��u�u�0�1�>�f�Wϻ�Ӗ��P��dךU����&�2�u�"�-��ԜY���F��V�� ���1�9�n�0�3��;��