-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B+��y���߇x��!�:�m��Ϝ���ƴF��^	�����'�?�6�o���(��L���"��RT��Dʟ�;�4�,�g�f�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�CחX���|�g�d�u�8�$����Y����\��'�����0�!�u�:�'�/����s����_
��^	��ʇ�&�'�0�_�z������ƅ�@��Z��ʜ�!�'�4�u�9�2�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�x��%�2��������\��Y��U���9�8�;�&�6�0�����˭�P��[��Yʡ�u�0� �0�w�3��ԑT����z4��^��ʢ�!�u�-�:�2�>�������g�������;�u�;�9�3�.��������Z��YחX���8�8�'�u�1�/�9Ͻ������
��ʸ�8�'�u�3�%�����Y����@O�V �������m�_�z�}�$�������(��V��ʴ�0�g�4�1�d�}�9������P
��\N��U���u�0�0�<�w�4��ԑT���	��^ ������0�3�6�2�)�M��Y�Ƙ�Z��X�����u�!�'�&��>��������@F��T������u�&�0�'�>��������[ǶN�����0�u�0�0�w�2�����ƻ�_
��D��ʴ�6�0�3�6�2�)����Ӊ��@%��Q*��Y���u�u�=�u�2�4��������\��YN�����1�'�u�;�w�2��������p	��`�����=�2�{�x�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���lǶd�U���0��<�=�6�9��������[F��[�� ���'�u�m�7�#�W�Z��Y����r$��-��;���u��u��2�
��������w��`�����u�u�0�1�:�1����Y����A��C�� ���'�u�<�0�w�<���Y�Ɓ�JF��Y��ʦ�'�4�<�0�6�.����Y����F��	��U���=�7�!�u�>�)�ϩ��ƭ�@
��RחX���u�1�!�u�6�8�Z�Զ����A��R�����&�u�0�0�$�9��������H��[UךU���u�0�0�;�:�/����݇��lǶN�����&�&�!�4�$�<��������A��6�����:�0�<�n�;�?����,����~]��D��;�����:�%�9�3����5�����C�����'�;�9�!��3�}������v��T �����_�0�0�<��}����
����[��N��U���7�:�0�;�m�}����B����u��C'�����u�u�u�;�5�2����C�ƪ�_��=N��6����1�=�u�w�}�W�������V��V ��U��!�u�m�o�w�e�}���=����Z��N��U��<�u�;�0�2�}����Y����\F��T��D��u�>�#�'�;�>�W���Y����]F��C��ʧ�;�0�g�!�w�}�J��P���A�N������>�-�u�w�g��������T��=d�����0��1�u�w�}�MϷ�Y����_	��T1�����}�u�:�;�8�m�L���
����U1��N��U���u�;�&�1�;�:��ԜY����V ��C��U���o�<�u�!��2����������R�����d�1�"�!�w�t�}���
����Z��X��U��<�u�!�
�8�4�L�ԜY����G��N��U���o�<�u�!��2����������C�����d�1�"�!�w�t�}���
����|��N��U��:�!�&�1�;�:��������X"��V9�����u�:�;�:�g�f�Wϭ�=����R
��~ ��U���;�&�1�9�0�>�}���
����e��S!��U��:�!�&�1�;�:��ԜY����G��~ ��U���o�<�u�!��2���Yӕ��R��R!��U���u�u� �u�#�����B����@'��E��<���u�u�u�;�$�9��������G	��N�����u�|�_�u�$�9����6���F��X�����9�2�6�#�4�2�_�������V�S�����'�h�r�r�l�}��������F�N��U���&�1�9�2�4�+����Q����\��XN�N���&��0��#�}�W���CӉ����h�����0�!�'�a�w�2����I��ƹ��T��:���u�u�u�u�"�}��������E��X��Bʱ�"�!�u�|�]�}��������Z��CN����&�1�9�2�4�t�}���Y����P(��=d�����!�6� �0����������KF��=d��Xǣ�:�>�&�2�#�/�}���T����X9��P�����6�;�!�;�w�����Y���F���*���<�
�0�!�%�j��������\������k�e�|�_�w�.����Y����Z��Y-�����u�u�!�
�8�4�W��^����9F��^	��ʦ��8�1�'�w�}�W���Y����_	��T1�����}�u�:�;�8�m�W��Q����A�^��N�ߊu�<�;�9�$�����6����_F�N�����2�6�o�u�g�f�Wϭ�����@��S������9�u�u�#�����&����\�
�����e�u�h�}�#�8����I����F��P ��U���4�4� ��;�}�W��
����\��h�����>�4�4�<�#�p�W������F��F�����h�r�r�n�w�.����Y����V ��s��U���u�u�!�
�8�4�(�������p	��`����1�"�!�u�~�g�WǱ�����A��UךU���;�9�&��#��������	F��S1�����#�6�:�}�w�2����I����N��_��H��r�n�_�u�z�6�����ơ�K9��Y��U���=�9�u�<�?�)����s�ƭ�G��B�����u�u�!�<�0�W�W�������VF��R��ʦ��<�0�;�8�?�W���Y����Z��[N��Uȡ� �w�_�u�6�)����Ӌ��l ��X��U���<�2�_�u�#�/����Y����U��B��ʦ��<�0�;�8�?�Mϭ�����Z�V�����0�<�_�u�z�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��ƹK�D�����9�1�;�u�z�W�W��1����Z��_�����3�'�1�!�w�<���Y����[��Y��U���4�<�;�!�!�1������ƹK�S��ʢ�<�0�<�u�8�)�Ϻ��ơ�^	����U���!�!�0���?����Yӯ��@F����U���u�0�u�=�w�2����������GN�����2�u�<�6�w�5�Ϭ�	����V��NN������>�_�u�z�}�Z����ƪ�A��z/�����4�=�&�2�2�)���� �ƨ�G��V��U����d�6�6�2�}����Ӓ��l�C�����4�0�:�,�w�(�W���Y����	��C��8���u�,�:�9�w�}����W�Ƙ�Z��X��U���u�u�x�u�%�-��������J	��[��U���!�0�3�:�w�;����
����_��X�����6�4�;�:�w���ԜY��ƹK�d��ʰ�1� �u�<�?�)��������\ ��D*�����<�u�<�;�;�q����Y����R
��Y��U���u�<�=�!�2�>�����ƿ�w�������{�u�=�&�>�}��������Q��B�����=�u�u�x�w�<����Y����V��_�����<�0�:�6�%�u�����Ƹ�VF��gZ�U���0�:�!�<�2�q�W��Y����J	��Y��U���1�&�7�0�#�8�1���Y������
��ʲ�<�2�!�u�?�0�������K��V��[���:�u�=�&�%�<����Y����@��C�����>�0�4�9�$�2�W���Y����E��VךU����r�u�;�>�8����=����F����ʢ�u�:�9�u�%�-����	����Z��C��ʴ�u�0�9�_�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l�C��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�x�w�<�ϓ�����F�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�u�x��}����Y���� �������u��9�,�6�>����Ӏ����C�����9�"�0�u�2�3����Y���w��a�����4�0�6�0�#�9�}�������] ��=N�����&�}�4�%�2�1�9���Yӄ��ZǻN��ʧ�&�;�
�1�2�����:����F��R ךU���u�&�'�!������Dӕ��R��R'�����&��!��;�9��ԜY�Ʃ�WF��d�����%�:�0�&� �4������ƹK�d<�����u�0�:�,�w�
�����Ƹ�VF��C�����,�"�0�u�!�/����Y����R
�������x�!�0�&��)� ���Y����VF��V��U���0�<�u�<�?�}�6��� �ƾ�R��E�����8�8�'�u�w�p�W���Ӓ����S
�����{�_�u�x�?�2�(�������~��EךU���=�:�
�u�$�<����Y����G��C=�����x�=�:�
�w�.����<�ƿ�d��R+�����u�x�#�:�<�<����������S
�����_�u�$�4�6�8����CӃ��Z��@��[���4�4�0�:�.�u�#���Y����V��^�����_�u�u�u��)� ������X"��V9�����u�x�<�u�>�)����Y����\��Z��]���u�u��8�;�����D�Ɵ�^��t�����u�x�u�;�w�)�(������F�D�����u�u�h�u�$�<����Y���F���U���
�:�<�
�2�)�ǵ�����W��N�����u�|�u�u�w�.� ������[�D�����;�:�7�u�z�}��������T��N��Uʦ��1�0�&�w�`�W�������@/��N��X���;�u�!�
�8�4�(��������Y��E�ߊu�u�u�&�6�<����Y����@"��V!��&���n�u�x�:�#�.��������V��EF�����<�!�x�u�8�3���s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���u�x�u�4�6�<�Ͻ�������Y	��ʡ�0���m�w�p�W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l�C�����:�!�:�u�>�8�W���Y����_��SN��U���!�u�4�6�w�5�W���������VךU���:�u�=�u�4�(�����Ư�R��=N�����1��;�'�;�g�WϮ�����5��G�����|�u�7�2�9�}�WϷ�Y����]��S	��&���9��>�-�w�5��ԜY���K��E��U���7�0�u�u�w�.�3���.������S�����4�0�;�_�w�}�W��Y����V��N��Uʦ��1�0�&�"����Y����W��D'�����u�u�x�u�6�<�!������F�N��U���&�<�u�=�w�4����8�ƥ��������y�1�9�,��)�!���ӄ��R��O�����u�u�x��4�>����Ӆ��C��V�����!�0�%�%�;�3�W����ƣ���+�����0�:�,�u�w�}�Z���+���g����R���0�1�1�<�w�5�W���Ӊ��G��z/��Yʷ�6� �0�!�2�9��ԜY���K��[��U���;�!�0�6�6�3��������F��D�����%�%�9�;�3�>����Y����R��=N��U���x�#�9�1�#�}����Y����w5��I�����'�4�u��$�}�W����Ƨ�Z��~ ��ʡ�0�_�u�u�w�}��������W"��R�����!��9�1�;�u�W������F�D�����9�1�;�_�w�}�W������F������4�<��,�k�}��������W"��Y�����:�>�#�'�;�>�^���s���F�N��U���u�u�u�u�w�.�3���/����z������>�#�'�9�4�p�W������]ǻN��U���u�3�_�u�w�}�Wϻ�ӏ��9F��Y
�����&�u�4�6�3�������ƓF�>��ʴ�:�2�:�!�"�.�����Ƣ�K��v-��ʡ�0�6�4�;�w�.�3���.����F�R�����!���!�4�f�Wϭ�8����@��CN��U��&��1�0�$�(�;���s�ƿ�w��x��U���u�i�u�&�6�<�������@��C����� �u�i�u�$�<����������R�����n�u�&��4�0����6���F��s��#���1�9�}��2�>����L��Ɠ9F�N�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�u�x��8��������r+ǻC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u��)����
��ƹ��T��]���%�0�9��~�}���������E�����1�0��8�;�����Y����9F�N��ʦ��4�<�2�8�;�J��Y����9F�N��U���4��1�u�j�.�4���8����9F�N�����u�u�u�u�$��������@��[�����6�:�}�&�3�/����P���F�R ����u�u�0�1�>�f�Wϻ�Ӗ��P��=��4���0�&�_�u�z�}����Y����]��O��U���9�u�3�1�;�$����
����W�������1�!�_�u�z�.�6�������V����ʱ�'�6�9�u�8�}��������~��E��U���6�u�<�9�:�6�}���TӒ����Q�����&�7�u�;�w�$����������
������<�u�&�6�>����Ӏ��9F�N��U���0�!�4��w�3��������C�������!�0���o�l�������9F������u�$�:�3�2�2����<����U+��X��Oʰ�!�!�u�:�<��4���4����JF��c"��U���2�;�'�6�:�-�_���Y����p	��`����u��0��3�5�W��Y���Z��P��U���%�'�u�4�w�W�W���Y����_��\ ��H���4�%�0�9��q�W������G��X	�����u�u�&�:�1�<����Gӕ��\��V��U���x�<�u�&�3�1��������AN��X�����x�u�:�;�8�m�}���Y�ƿ�p	��`��U��u�&�:�3�2�}�W���Tӏ����h���ߊu�u�u�&�6�����Y����@4��v
��Y���u�x�<�u�$�9��������G	��N�����u�|�u�u�w�.�4���-����[�D������%�n�x�w�(�W���&����P9��T��]���0��1�=�f�9� ���Y��ƓF�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�x�u��i�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�dךU���=�:�
�u�&�.�C�ԜY�˺�\	��VN����� �4�:�u�6�.�}���T����X9��t��&���9��>�-�w�p��������rF��s��:���'�_�u�x�?�2�(���<����@��C�����9�}��0�4�2���s���E��\1�����g�&��!��1����Q����A��T��\���x�#�:�>�6�>�W�������w��N����>�4�6�6�9�.�6�����ƹK��_��*�����&��#������Χ�E��[��^���u�x�#�:�<�<�����ƿ�r��Z!�����x�=�:�
�w��8�������F�A�����6�u�&�'�0�(�}���T����X9��T+��U���4�4�4�<��$��������XM��=N��X���:�
�u��4�0����Y���F��s��M��0�!�!�u�8�6�2���	���a2��=N��U���0�<�u�4�w�W�W���Y����@��t����u��'�!�9�5���Y����]F��X�����h�3�9�0�w�}�Wϵ�����_��EN��Kʳ�9�0�u�u�w�}�W��Y���Q	��R��O���4�&�_�u�w�2�ϳ�	��ƹF�-��U���u�u�u�k��0�������F�N��U���u�u�u�x�w�3�W���&����Pl�N�����u�u�u�u�j�}��������A
�N��U���u�u�u�u�w�p����
����\��h�����d�u�:�;�8�m�}���Y�Ư�]'��N��U��u�&�4�4�6�4�3�������P
��\E�Y���x�<�u�&�3�1����Y�����v\��U���u�k�&��#������Χ�E��[��^���u�x�u�;�w�)�(������F�T,��U���u�u�h�u�$�2����
���F�N��U���u�u�u�x�>�}��������l��C��D���:�;�:�e�]�}�W���<���F�N��U���4�4�4�<��$��������XM��N��Xʼ�u�&�1�9�0�>�W���YӅ��F�N��U��&��0��#�}�W���Y���F�N��U���u� �u�!��2��������R��S�����|�u�u�u�4�3�W���Y���F��s��#���1�9�}��2�>����M���K��YN�����:�<�_�u�w�}�'���Y���F�������y�u�u�w�}�W���Y���F�N��Uʦ�1�9�2�6�!�>����Nӂ��]��GךU���u���!�w�}�W���
����F��CB��U���u�u�u�u�w�}�W��Y����@��[�����6�:�}�b�3�*����P���F��v�����u�u�k�:�2�q�W���Y���F�N��U���u�u�x�u�"�}��������E��X��Lʱ�"�!�u�|�w�}�WϽ�����_��S�R��n�u�u�u�w�}�W���Y���F�N�U���u�!�
�:�>�W�}���Y����9