-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B/��B�����;�f�6�#�3�p�W�������w��u�����u�'�2�;�;������Ɯ�z��Z������!�o�d�w�<����Y����9K��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�w�>�W��Jӥ��J��_�����;�9��&�%�0����:����A��X חXʔ�9��2�!�w�8�������}��X ��U���!� �0�!�w�3����ӯ��\��C�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z��Y����\��=C�Uʁ�<�u�:�%�9�3�W�������G��^ ��ʦ�8�9�;�{�w�2�W���Ӕ��\��RN�����4�<�;�x�w�}��������F��R�����#�'�<�;�w�;����Y����\��CN��ʾ�#�'�9�6�]�p�Wϻ�����F��SN�Uʚ�=�'�#�9�2�}�����ƿ�C��C�����=�&�!�8�y�p�}��YӲ��@F��Z�����!�>�&�<�w�����Y����@"��V8�����y�4�1�%�8�(��ԑT����@"��V=�����y�&��!��1����	�����������<�{�u�&�6�<�����ƭ�G��[חX���6�8�&�<�w�*�W�������@"��V(�����8�9�1�4�3�.�3���*����W5��G��[���=�_�x�u�u�4�����Ƹ�VF��X��U���2�0�0�!�w�3�W���Yѕ��\�������,�1�7�u�9�W�Z�������R
��V�����u�,�9�{�w�5�����ƹ�V��V��U�����7��#�/��������[ǶN��8����4�;�!�2�9�����Ʃ�R��DN�����9�u�9�2�2�q����Ӊ��D��_N��ʳ�9�0�_�x�w�4�W���s��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�_�<�'�%�}����s�ƹ�VF��R�����:�<�
�d�c�<��ԜY����Z�� �����
�!�{�9�l�W�����ƻ�A��N��ʢ�'�{�>��y�1�L�������\��g�����9�!�0��'�<��Զ����JF��~ �����%�<�2�:�w�.�������F��V�����u�u�u�u�w�g��������AF��Y	��D���:�d�u�h�f�f�Wϵ�	���F�N��U���u�u�;�<�#�:�Ϭ������X��O���u�n�%�'��}�$�������}�N��U���u�;�&�1�;�:��ԶYӕ��\��a��U���u�u�u�u�9���������9l�D*�����<��u�u�w�}�MϷ�Y����_	��TUךU���!��u�u�w�}�W���Y�ƥ�5��s��*����6�d�1� �)�W���s�ƿ�w��q�����%�0�u�o�8�)�$���������TC����!�u�|�o�w�2����D�Σ�[��
P��R���_�u�&�4�6�8��������WF��X��&���4�4�!�>�'�p�W������F��F�����h�}�!�0�$�c�G���B����@"��V8�����8�9�1�u�w�(�W���&����P9��T��]���6�d�1�"�#�}�^��Yۉ��V��	I�\�ߊu�&�0�=�>�}�W���Y���	F��CN�����2�6�o�u�g�}�L��ӣ��]��d�����f�6�_�_�%�5��������g*��QN��<���!�4�%�<�0�2�W���s���E��\1�����'�_�u�x�?�2�(�����ƓF��Y������0�6�:�<�}�W������V��V ��U���:�f�o�u�l�W�W��������V�����4�&�0�<�;�9���� ����\F��D��U���,�!�0� �2�}������ƹK�^ �� ���u�;�!�0�u�8��������F��N��R���<�0�,�&�6�1�Ϫ��Ƹ�VF��E�����x��6�4�6�)����W����J��N�����4�4�'�4��}�Ͽ����X5��_�����:�e�u�3�$�9��������G	��\*�����!�x�u�:�9�2�G��Yӕ��]��D�����0�u�u�u�w�}����=����A��h��H���!�0�&�k�8�5���^���lǻ�����&��!��;�9����Y�ƿ�W9��P�����:�}��6�f�9� ���Y���F��C����e�|�_�u�$�:����
����u��CN��U���u�8�9��#��������	��R��Kº�=�'�h�r�p�t�}���������V�����1�u�u�o��<��������J9��S�����'�h�}�!�2�.�I��P��ƓF��P ��U���4�4�0�4�2�}�W��*����w��v�����o�u�:�=�%�`�_������V�UװUʦ�2�4�u�&�2�5�������\��C
�����u�h�r�r�]�}�����ƿ�p	��C8��0���9�u�u�:�;�<�!����Χ�C�
�����e�u�h�}�#�8��������lǻC�>���u�;�!�0��.��������Z�C�����u�=�8�7�>�:�����ƻ�G��_�����_�u�x���)����
����[��D��U���4�}�;�!�2��W������F��C�� ���>�0�u�u�#�4��ԜY����Z��RN�����3�&��!��8�W���Y���	F��P ��U���w�'�0�n�w�<��������V��X�����4�4�<��2�}�W��
����_F��L�� ���_�u�!�'�5�)�W���	Ӊ��@��B ����� �9�u�u�w�4��������A��d�����<� �0�>�2�}�ϭ�.����Z��[N��U���o�&�2�4�w�.�U�����ƹ��E�����0�%�:�u�$�<����
���F�T�����9�<�u�!�"��}�������F��\��U���&��!��4�3�W���Y����@��V�����'�0�n�_�w�p�#�������@F����U���
�4�:�!�w�8�Ϻ�����]��R�����;�4�9�y�5�}�������K��_�����4�9�;�u�>�4�Ϭ�	����9F��C�����u�4�
�4�8�)�W�������F��C�� ���8�-�3�;�"�}�ϭ�.����Z��[N����4�u�&�w�u�W�W�������VF��O1�����u�3�&��#�����Y�ƿ�T����W���_�u�!�'�5�)�W���&����F��QN��1����6�;�u�w�4�������]Ǒ=d�����_�u�x�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��Y���z��CN�����;�_�u�x�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F��R�����u�0� �'�3�<��������UF��s��<���&��!��;�9����
����R��G�U���u�;�u�&�3�/����Q����@F��R�����0�;�u�4�$�9�����Ƹ�Z��X�����u�;�_�u�z�4�����Ʃ�@��^�����&��!��w�5�����Ơ�]��B�����&��1��6�3�G��U���F��s��#���1�;�&�:�;�}�����ƥ���X �����9�y�4�1�$�
�4������@��[
ךU���%�0�0�1�>�}�Ͽ�������G��Uʁ�<�u�&�&�:�1�Ϫ�Y������@ �����x�u�<� �2�h�EϷ�Y����k��Y�����-�a���"�8�W�������TV����U���%�'�:�6�~�W�W������[��[�����u�&�&�4�0�/�Ϻ�Ӓ��u ��C��U���0�7�0�u�3�8�W�������RǻC����8�'�#�u�>�4��ԜY��ƹK��N�U���;�>�#�'�;�>�J�ԜY���F�N��U���u�u�u�
�w�}�(���Yӹ��F��hN��U���u�u�
�u�w��W���&���l9ǻC�&���9��>�f�w�}�(���Y����F��h��	���u�)�
�u�+��WϢ�&����l9����	���
�_�u�x�w�p�W�������R��G��Uʩ�u�u�)�u�w�!�W��������N��U��u�u�g�u�w�m�W���H�ư�F�N��U���u�u�u�u�w��(���&ӹ��l9��h1��*���
�u�
�
���(���&����l9��h1��*���u�x�u�&�6�<����
���lF��h1��	���
�
�u�u���(���&����lF�h1��*���
�
�
�
���W��Y���F�N��U���
�
�
�
���(���&����F�N��U���u�u�u�
���(���&����l9ǻC����!��9�1�9�}�W���Y���F�N��U���
�
�
�
���(���&���K�N��U���u�u�u�u��}�W���Y���9��h1��U���u�u�u�u���W���Y���F�h1��*���x�u�&�0�?�4�_���Y���O9��h1��*���)�u�u�)���(���&���F��h1��*���
�
�_�u�z�}�Z���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǑN�������8�<�m�}��������R��R-��;���u�7�2�;�w�}��������l��RF������>�-�u�?�3�}���Y�ƪ�AF��^ ��U���>�%�x�u�8�-�W���Y���F��R��U����#�'�<�9�2�W���
Ӊ����[�����u�:�u�<�>�:�W���Y����@%��Y�����4�d��u�j�.�4�������zO�^�����u�u�u�x�w�5����?�Ƹ�R��R�����!�0�d�u�8�<�Ϫ�Y����}��X������0�0�4�2�}�W���Y���X��DN��U���8�!�u�;�"�8����Y����GF��CN�����u�<�=�1�'�4����Y��ƹF�N��Xʺ�=�'���w�3��������bHǻN��U���3�&�� �#�8�2����΅���Yd��U���u�u�&��#�����Pۍ��G��S��Dʱ�"�!�u�|�k�}�3���0�΅���C�����d�1�"�!�w�t�}���Y���F��s��#���1�3�'��w�`��������W/��=N��U���u�;�u�3�]�}�W���Y���}�������,�!�0�1�#�}���*����V%�������!�>�;�u�9�2������ƹF�N��Xʡ�0�1�!�#�;�9�������g���� ���u�:�u�=�w�.����[Ӊ��C��=N��U���u�3�&��#���������[�N��ʦ�� �!�0��(����PӒ��]l�N��U���&��!��;�$�Ǘ�Y����@"��V6���n�u�u�u�w�8�Ϸ�B���F�R �����n�_�u�u�w�.��������[��D*�����'�_�u�u�w�.��������Z�D�����9�,�1�_�w�}�W��Y����R��YN��ʶ�6�0�7�3�%�}��������F�N��U���:�;��6�g�`�8�������U��_��U���u�u�&���<����Y���A��R��U���0�=�<��;�a�W��B���F��Y
���ߠu�u�0�1�>�f�Z�������l��Rd�����%�:�0�&��.�#���=����]]Ǒ=N��Xʜ�%�!�&�8�;�3�W���Y������_N�����!�4�u�0�2�7�����ƾ�T��D��Yʡ�u�0�&�'�]�}�Zϩ�Y�����\��Wʴ�,�0�!�4��z�Y�������AF��RN��&���<�!�'�<�'�)�W���s�����Y	�����%��!�
�w�$��������W	��YI�����u��!��3�5�Wύ�Y����I��Xd��X���4�6�u�=�#�}�#���Ӄ��A������7�u�%�<�>�8�W���Y����\��[�����_�u��&�-���������C��R�����!��'�!�]�}����s���@��C�����4�%�0�u�j�u����
����G��DS�E���n�u�u�3�%�����Y����`��N���ߊu�u�u�&�6�<����*����V��F�����<�!�x�u�8�3���Y����@"��V(�����|�_�u�u�9�}����s�Ʃ�WF��X��ʇ�&�/��!��/��ԶYӴ��Z��V�����1�u�'�6�$�u��������]�N�����u�u�&��#�����*����V�
N�����&�k�:�=�%�`�P���P���F��EN�����u�:�>�%�z�}����Y�����V�����1�4�%�0��t��������[K��S�����|�i�u�&�6�<����ۯ�9F���U���%�_�u�;�w�/����Y����I��C�����n�_�u�&� �����E�ƿ�d��V����u�&��!��1����	����[��D*�����<��0�n�]�}�Zϛ�Ӊ��z��CN�����;�_�u�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s���WF��{U�