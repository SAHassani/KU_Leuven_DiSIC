-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:��:�>�!�9�Z�������	F��_ �����8�;�x�u�%�:����)����P��g6��*��`�_�x��#�g�F������W��CחX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�_���K����p	��E��ʛ�!�:�4�u�9�)�����Ə�A��V�����u�9�u�<�?�.�%�������K��V������&�'�8�9�.�>�������z��E�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s����F��D�U���&�3�9�u�%�<�����Ƽ�\��D��U���6�u�:�u�?�}��������9K�N��U���u�<�!�'�8�<���Y����[��DN�����0�u��8�%�>��������@l�N��U���u�u�'�6��)��������GF��X��[���_�x�u�u�w�}�Wϊ��ơ�W�������4�;�"�6�;�(����Ӄ��A��^�����'��9��w�.����s���F�N��U���0�u�;�&�?�.�W���Y����R4��S/������3�0��{�4�W���Ӓ��]F��[�����!�0�x�u�w�}�W���Y����V��B��ʦ�6� ��!�x�}�����ƺ�_��@��U���6�8� ��;�9�������K�N��U���u��4�0�$�2����Ӑ��Z��E�����8�8�;�u��<��������@��C�����0�4�;�x�w�}�W���Y�ƺ�_��Q��R���0�6�:�>�6�)���� ����l�=C�U���u�u�u�&�6�<����0�ƥ�W��C�����=�'�u�&�9�*����Y����VF��D��U���:�!�0�8�:�/��ԑT���F�N��Uʓ�'�>�4�%�2��������J��s��'����1�0�&�1�.��������Z��V �����0�_�x�u�w�}�W�������GF��R
��ʼ�;�'�u�=�w�4��������@F����U���3�u�0�<�#�/�Lϊ��ƥ�9K�N��U���u�;�0�0�w�8����Y����w�������;�2�:�%�w�;����	����V��T��U���6�u�0�;�]�p�W���Y�����E�����6�;�7�u�"�5�Ϫ�Y����^��E��Yʰ�0�u�=�;�>�}�ϰ�ӟ����S�����x�u�u�u�w�}�W���Y����V��T�� ���<�;�u�4�>�}�3���+����W��D������u�4� �$�<����I���W�C��U���u�u�u�;�w�l�U�ԑT���F�N��U��x�u�&�u�?�}����ӂ��RH�r�����d�:�u�=�w�<�Ϩ�����R��=C�U���u�u�u�u�w�}�WϷ�����]��R�����"�0�u��#��!���Ӈ��V��@חX���u�u�u�u�w�m�W���,����[��R��ʻ�"�&�u�4�6�}�2������	��C�����u�4�<�u�6�<�}��Y���F�N��U���u�;�9�1�9�}��������[��D*�����4�<�u�&�2�)�^�ԑT���F�N��U��x�u�&�u�?�}����Y����@��V�����u�u�u�u�w�}�F���GӲ��@F�� ��U���4�<�u�3�$�)�}��Y���F�:��ʦ�2�4�u�&�#�0�W�������G	��s��#���1�;�_�x�z�}�W���Y���z��V��U���,�9�&�}��8��������w��NG��ʶ�9� �4�0�#�8��������]��C��U���u�u�u�3�2�}�$�������z��D������<�u�0�9�}��������C	��^ �����u�:�u�=�]�p�W���Y�����T�����u�0�1�u�8�/��������r%��Y��Mʶ�:�>�u�,�;�.�������F�N��Uʦ�!�'��9��}��������GF��\��Gʶ�6�0�u�:�1�:�����Ƹ�VF��P�����_�x�u�u�w�}�Wϳ�����A�������u�9�&�d�4�>�Ϫ�Y�������� ���1�!�u�'�:�0����U���F�N��Uʓ�'�!�<�u�2�.�ϭ�����e��SN��ʦ�4�4�0�1�3�/��������]F��RN�����1�x�u�u�w�}�W���Yۍ��G��[�����|�6�6�0�w�3����Y����_�CחX���u�u�u�u��}����Y����P��R��ʢ�<�0�4�1�#�8�W���ӂ��RF��X������u�4�4��0����U���F�N��Uʁ�u�4�6�u�?�}�4�������c��s��ʢ�u� �!�=�!�}����Y������D*�����<�0�z�_�z�}�W���Y�����T�����0�u�3�0�w�����������R��U���u�;�u�9�4�}����Y����Al�N��U���u�u��!��1����Y����c��b ��ʢ�9�u�0�4�w�5�W�������Z����U���9�u�:�6�2�)�}��Y���F���U���:�,�"�<�2�.����Uӕ��G�������<�0�4�<�9�9� ���Y����R/��^��Z���x�_�x�u�w�}�W���-����Z��^ �����,�!�'� �?�)����������^�����&�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��Ɠ_��V�����y�"�'�n�w�(�Ϸ��ȿ�W9��P��D��{�9�n�u�"�8����W����A��D�����_�u�&�u�8�6�'�������Z��D*��[���n�u� �0� �/�Y���?����z��E����u� �0�"�%�s����	݇��l��Y��ʓ�4�!�;�0�'�/�����ƥ�9F��R �����u�u�>�4�'�8�'��� ����	F�������u�4�2�u�w�2�E��Y��ƹF��x�����>�4�!�'�m�4�W�������A��RN����u�h�f�_�w�}�9�������@��b ����<�u�4� �6�}�J��P���C	��d��Uʆ�8�9��>�m�4�W���&����P]ǑN��X���#�'�u�<�2�.����:����R��E��U���0�u�<�!�%�4�W�������V��V��U���&�=�&�{�w�}��������PF��^ �����4�n�u�u�$�5����Cӏ��c��R1�����%�0��'�.�1�Z�������V�C� ��m�_�u�u��)�>��������U�����_�u�u��#���������| ��R��U���;� �&�2�2�o����&�Χ�R��R�����9�x�u�:�9�2�G��T�ƙ�TǻN��1�����%��m�4�W������F��@ ��U���u�x��m�f�}�Wϭ�����c��fN����<�;�1�d�w�2����I���F��@����u��6�8�"�����CӉ����[��N���u�&�6� ��)�W����ƈ�G��C1�����%�0��'�.�1�Z�������V�N�U��{�_�u�u��>����(����F��V�� ���}��8�9�$�8�4�������\��XN�\���x�u�a�{�]�3�W�������V��E�����n�_�'�=�#�>����+����UF��V�����%�'�6�9�4�}��ԜY����6��D�����<�u�'�4������
����J��_�����:�e�u�3��<��������A	��D�����!�u�:�;�8�m�L�������w��v��ʼ�u�'�4�}�6�(��������X�X�����;�1��'�.�)����)����@��P;�����:�;�:�e�l�}����Y����V��v��ʼ�u�'�4�}�9�)��������Z�N��U���;�1�a�u�8�3���B����J��v�����
�u�&�4�%�$����	����V��T��Dʱ�"�!�u�|�8�}�����ލ�J9��\ ��%���0�&�;� �>�.��������l�C��U���9�4��!�>��W���������Z������6�0�d�3�*����PӉ��q	��R�����'�>� ��8�8����,������Y��E��u�x�u�9�w�5�W�������a	�������=�u�4�0�3�)�W�������F��D�����=�<�u�3�3�)�W�������A��N�U���%�:�4�4�2�.����������C�����u��!���-�>���Y����VF��[N�����<�;�9�4�$�:����
���F��RN�����;�<�0�4�0�3����Y����V��CB��ʶ�0�!�u�u�"�)�Ϫ�	�Ƹ���G��ʡ�0�%�'�_�w�p��������G�x ��U���8�;�u�u�9�.����������B��U���1�<�0�!�2�9��������9F��N��<���!��,�!�>�}����QӍ��^��D>��6���0�x�d�1� �)�W���Y����Z��S_�����
�}��8�%�>��������@F��@ ��U���_�u�x�u�%�<�Ϸ�����W��RN�����&�!�u�<�2�4�Ϫ�Ӆ��G�������u�;�u�4�4�}��������A��^�����u�;�!�0��2�"���
���@��V��1�����9�1�>�8�MϜ�����e��X��1����9�1�0�6�}�W�������V�S�����'�u�k�3�;�8�L���
����_F��E�����o��4��.�)��������W"��V��Dʱ�"�!�u�|�m�}�������N��_��U��}�!�0�&�j�}�G���P��ƹ��Y�����'��9��.�g�5�������G��h�Uʦ�2�4�u��6�8����Y����V'��h�Uʦ�2�4�u��#��6�������A�*�����
�}��8�;�.���������Y��E��u�&�2�4�w���������JF��u�����4�'�-�!�]�}����ӕ��G��N'��U���4�4�'�
�l�}�����ƿ�R��E��Oʜ��!��,�#�W�W�������r��Z8�����,�o��:�2�3��������F��P ��U���6�8�'��m���������9F��^	��ʦ�6� ��,�w�}����8����l�D������6�8� ��$�W�������A��d�����4�u��6�:�(�6���Y�ƍ�P��E��N�ߊu�x�=�:��4���������X�����1�_�0�<�]�}�Z���������R�����0�&�:�u�1�.��������WF�������=�u�<�0�>�8��������]��YN��ʅ�:� �<�&�]�}����
�Ο�^��t�����0�<�_�u�w�;��������T��V�����|�!�0�_�w�}�W�������R
��g��U��&�4�4�;�6�4�'���Q����R/��V��%���r�<�=�x�w�2����I���@"��V'�����n�u�u�0�3�4�L�������A	��D����u�x��0�1�/�Ϯ�����Z��B ��U���0�u��!����������V��NN�����4�<��9�.�>����W���K�y��Oʦ�4�4�;�4�>������ƿ�R��Y>�����u�'�u�:�w�4�Ͽ�����l�N�����4�<��,�g�u�^��Y����R/��V��%���}��!���1����Ԏ��[O��N��X����!���'�}�Ϻ�������N�����>�6�6�0�w�3����5�ƨ�R��Z@�����8�!�=�&�#�8�'���,����F�C�����'�8�;�y� �}��������Z��^��ʡ�0�3�'�!�'�2�����ƹ�Z�N�����4�'��e��t�K���=����]6��R'�U���&�4�4�'��m�_���E�ƿ�R��Y>����_�u�0�0�6�8��������D��N��ʆ�6�;�0�u�9�6��������p��RC����!�u�u�0�2�<����Y���z��^�����=�u�<�&�w�1����Y����[��E��U���3�0�u�=�w�4��������@����ʺ�_�u�u�x�2�>�W���Y����D����U���u�0�0�u�>�3�����Ư�V��V�����!�'�6�'�>�.�}���Y����@��NF�����0�|�e�u�j�.����Q����]��UךU����4�!�4�4�/�_���0����N��R�����'��9�n�w�}��������zN��T'�����e�u�h�}�#�8���Y���l�N������,�}�%��9����P���	��R��H���e�|�_�u�w�p�W����ƿ�R��R�����&��3�0��}�ϳ��Ƹ�VF��X�����<�0�<�0�3�1�Ϭ�����^��D@ךU���'�6�&�}�6�-����P�����^ ךU���u�3�'�&�9�����*����V%��N���ߊu�u�u�u��<�'���Q����]��F��1����9�1�0�6�}�W�������V�S��1����%�}�%��9��������e��S*�����u�u�:�;�8�m�W���=����V��S
�����3�0��}�'�����B���F��Y
���ߊu�u�;�u�%�>���Y���F��R ��&���9�&�0��4�8����Y����w��<��ʔ�1�0�&��1�8�W�������@F��=N��U���!����1�8�6���*����W��^��I����4��%��-�>����Χ�R��V��1���,�x�d�u�?�3����	����V��T��H��0�&�u�:�?�/�W���^���9l�N�����!��:� �>�.�}���Y����ZF��_��ʾ� ��:�0�$�3�"���
Ӂ��V��Rd��U���x�#�:�>�2���������c��b �����u�u�x�=�8��W�������R��F��D�ߊu�u�u�x�?�2�(���*����p��~ ��&���!�4�6�'��-�>����Υ�OǻN��U���=�:�
�u��<����
����V'��=��<���-�}�x�|�w�}�W������l��s��'����1�0�&�1�.����
����a��x�����,��6�;�2�t���s���F�A�����&�!�'��;��ϭ�����R
��E�����1�-�}�|�w�}�W������l��g�����u��4�0�%�u�������ZOǻN��U���=�:�
�u��)�%���8����@��Q��:���&�4�4�1�3�;�����Ο�P/��R���ߊu�u�u�x�?�2�(���=����]0��^
��1����9�1�'��t���s���F�A�����&�4�4�;�>�8�W�������zN����\���u�u�x�#�8�6�ϭ�����c��fN�����'��e�}�z�t�W���Y����[	��h��1����!�4�<�w���������JN��T'�����<�_�u�u�w�p����&�ƿ�R��B�����4�'���4�3�������F�C�����4�&�4�4�"���������5��~ �����|�u�u�u�z�+����ӕ��P��Y'��4���8�'���4�3�������F�N����>�4�&�6�"��&ϭ�����A��d�����|�<�d�_�w�}�W�������RF��T��:���4�<�u��4�0����8����C��S��]���u�u�u�x�!�2����
����^)��{��U���6�8�'���>����Pۏ�F�N����>�4�&�6�"�����(ӕ��P��E��&���;�0�|�<�]�}�W���T����X9��D/�� ���!�u��6�:�(�6���Q����]��F�����u�u�x�=�8��W�������G7��v������,�}�%��9����P���F��E��<���'��:� �>�%�W�������\��q�����0�%�'�6�9�)�_���P���F�	�����u�4�u�_�w�}�W���Y����C
��g�����u�k�>�4�'�8�'��� ����F���U���0�0�u�4�0�}�W���K���l�N��U���>�#�'�9�4�����Y����|��T�����!�'�u�x�w�3�W�������A��RN����u�h�f�u�w�}�W�������]��Y��U���h�u�<�d�~�}�W���Y���K�^ �����2�'�o�u�]�}�W���Y������FךU���u�u�u�4�'�8����Y���F�N��U��u�4�%�0�;�q�W���Y���F�N��U���u�u�x�u�9�}�������F�N�����'��9��w�}�W���Y���[�D=�����9��,��4�3�������F�N��Xʼ�u�7�:�0�9�}�W���Y����c��R'��U���u�u�u�u�w�}�W���
����V'��=��<���-�}�x�|�w�}�W���Y����������_�u�u�u�w�}�$�������|��N��U���u�u�h�u��<��������`��Y
��\¼�y�u�u�u�w�p�W���Y����V��N��U���u�&�=�&��)�W���Y���F�N��Kʦ�=�&��,��>����Pۏ�F�N��U���u�x�:�!�"�.����Y���F�������9�1�u�w�}�W���Y�����C�����'�}�|�<�f�q�W���Y���F�C�����:�9�4�_�w�}�W���Y����R4��S/������3�0��w�`�W�������W)��D�����%��1�-��p�^���T�ƥ�F��D�����u�u�u�u�$�<��������F�N��U���u�k�&�4�6�/�>��Q����F�N��U���u�u�u�u�z�4�Wϭ�����9F�N��U����!���'��W���Y���F�
P��1����,�}�|�>�l�[���Y���F�N��U���u�;�u�<�9�9�}���Y���F��V�� ���9�1�u�u�w�}�W���D�ƿ�R��V��4����6�;�0�~�4�[���Y���K�X�����0�;�u�u�w�}�Wϭ�����R��S�����&�!� �u�i�.��������U��v��&���;�0�|�<�{�}�W������]��YךU���u�u�u��#�����Y���F�N��U��u��!��.�u�������ZO�N��U���u�u�x�u�"�}�������F�N�����4� ��u�w�}�W���Y���[�D*�������6�;�2�t���Y���F�N��Xʺ�!�&�2�0��}�W���Y����r��Z'��U���u�u�u�u�w�}�W���
����^'��~F�����0�|�<�d�{�}�W���Y����������_�u�u�u�w�}�6�������F�N��U���u�u�h�u��>����(۵��z��OG��X���u�u�u�u�w�p�W���Y����V�N��U���u�&�6� ��)����Y���F�N��Kʦ�6� ��,��-�>����Υ�F�N��U���u�x�:�!�$�:����Y���F������ ��9�u�w�}�W���Y�����T������6�;�0�~�4�[���Y���F�C�� ���<�;�1�_�w�}�W���Y����F��C8�����u�u�u�u�w�`�W�������_��E�����1�-�}�|�w�}�W���T�ƣ�GF��X�����u�u�u�u�$�>�������F�N��U���u�k�&�6�"�����0۵��z��OG��\���u�u�u�u�z�2�ϭ�����9F�N��U����6�8� ��}�W���Y���F�
P��4���8� ��,��-�>����Υ�]�N��U���u� �u�<�9�9�}���Y����T��E��U���0�4�0�'�4�3���s���@'��B�����%��1�-�w�`��������r��=��<���-�}��8�%�>��������@O�N�����u�|�_�u�w���������C��S��U��&�6� ��#�/�&Ǎ�����KO��y�����&�<�2�;�#�t�C�������V�=d��U���u�0�0�4�2���������P3��C<���ߠu�u�x��;�)�Ϯ�����Z��B ��U���&�=�#�u�?�}��������C��
�����u�u�x��w�8�ϱ��ƣ�VF��T��:���4�<�y�"�w�<�W���Y������@��U���u�=�u�<�$�}���Y�ƿ�P��x�����u�h�&�6�"�����������Z>�����<�2�;�!�~�W����+����