-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B5��P�����'�#�1�x�w�(����Y����q��Ed�U���2�;�9��8�8����!����R��=C�1���o�d�u�4�"�/�W��J���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�6�w�m�Dϝ�	����[��V������&�'�8�9�.�4�������\ǶN��ʇ�2�!�u�0�2�+���Y����\��'�����0�!�u�;�2�3�ϗ�����G��=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z�p�W���	����9K�N�����:�%�;�;�w�0���������������<�u��u�>�)����0�Ƥ�@F��R��X���u�0�0�<�$�W�Z���YӍ��V ��S��Xʦ�0�<�<�&�#�8� ���Ӊ��G��T�����0�!�{��;�}�Oϭ�	����V�C��U����!��1�?�p���������������3�!�0�1�#�}����
�ƃ�_�N�����!�1�_�x�w�}����	����W��N�����<�&�=�"�:�3�W������F��C�����0�!�:�u�?�}�������F�N��U���u�u�u��2�9����ӏ�� W�^ �����u�4�0�-����������Z��B�����u�u�u�u�w�}�W���YӒ����Y
��ʺ�0�4�<�;�>�}��������w5��@��"���u�m�7�!�z�}�W���Y���F�N�����&�4�1�4�d�}��������F��RN�����u�4�u�a�>�)��������K�N��U���u�u�u�u�6�9�F�������\��������0�3�4�#�2��������R��U�����u�u�u�u�w�}�W���Y����V�������u� �u�=�w�3����Y������SN��U���!� �6�!�3�p�W���Y���F�N��U���u�=�;�&�#�/�����ƀ�Q0��`@��,���6�;�>�0�w�-����NӉ��K�N��U���u�u�u�u�#�8�����Ʈ�G�N�����!�>�0�u�?�}�O�������Z��BחX���u�u�u�u�w�}�W�������]��_�����<�2�&�=�:�}�Ϫ�ӊ��GF��gZ�[���:�u�:�9�]�p�W���Y���F�N�����;�6�9�,�0�}����Y����Z����U���!�1�0�;�#�0��������K�N��U���u�u�u�u�1�/�F����ƥ�C��S��[���u�u�u��:�<����*�����E������6�&�2�2�)�W���Y����F�V �����u�4�_�x�w�}�W���Y���F�N����� �0�u��2�>��������Z��Y�����u�u�>�#�%�1����Y����Z ��DN��ʺ�0�6�:�>�9�}��������[��E�����u�3�x�u�w�}�W���Y���F��V������u� �!�5�}��������]��X�����0�9�u�u��8�������F�N��U���u�u�u�4�3�)�Ϫ�Ӆ��P��Z��U���%�4�0�4�>�3��������R�������u�u�u�u�w�}�W���YӅ��Z��Q��U���u�4�0���s�8���Y�ƭ�WF��D�����1�u��9�2�W�Z���Y���F�N��Uʲ�0�!�'�!�6�}�W���Y����R��NN�����u� �%�'�2�}��������9K�N��U���u�u�u�u�w�2�Ͻ�����F���� ���3�d�<�;�#�.�������@	�������x�u�u�u�w�}�W���Y����Z�������9�6�<�2�$�2��������VF��^��ʼ�u����]�p�W���Y���F�N�����6�9�{�u�z�}�W���*���F�C�����3�0�u�=�w�(�����Ƽ�A��R�����0�u�;� �w�3�W���	��ƴF�N��U���u�u�u�u�9�8��������p
��T������9�1�#�;�8�W���Y���F��V�D���x�_�x�u��8�������� ����ʳ�9�0�u�&�u�8�®�����_D�V �����0�,�&�8�;�/��ԑT����Z��RN�Gʼ�u�=�u�<�>�%�!�������w5��B��U���9�u� �e�d�-�������[F��YחX���8�1�3�6�#�2�϶��Ʈ�V��V
�����9�:�u�=�w�8����
Ӈ����X�����u�<�<�2�]�p�Z���Y������G�����4�1�0�u�?�}����Y����_��N�����!�;�u�'�:�)���Y�Ƀ�G	ǶN��G���'�4�&�u�9�}��������G	��C��U���!�%�0���?����ԕ��\F��R��U���x�u�u�<�0�8�1�������AH�v����� �&�4�0�d�}����YӲ����Y
��ʺ�6�'�_�x�w�4�W���Y����"��V��U���u�=�u�4�"�<�����Ƹ�VF��C��ʷ�!�u�<�9�5�}�Z���Y����_��^ ��#ʓ��{�x�_�z�}�#���ӈ��Q��X�����<�<�;�&�w�����
����V������>�#�'�9�4�W�Z��Y�Ƙ�VF��R�����!�u�=� �3�?�W�������@F��[���߇x�u�x�u�8�}�$���H�Ơ�R��_�����<�<�;�&�>�}�����ƣ�W����[��u�y�g�u�y�t�Z���Y����\��d��D���:�1�!�0�4�8��������D����&���&�0�u�<�2�}��������R��C��U���!�u�=�u�2�4����Y�����������=�u�;�{�z�}�W���?����K��[��ʾ�%�h�u�;�w�5����������Q�����&�u�&�u�?�.�������F�N��E���y�m�u�d�{�l�[��U����T��=C�U���u�u�y�`�w�q�W��Y���W�[�G���x�u�u�u�w�o�W��H���J�B��G���c�u�e�_�z�}�W���Y���F��N�Y��y�g�y�g�{�n�}��T���c��[��U���4�&�3�'�!�/��������T��C���߇x�u�x�u�w��[��Y����	F��A�����h�y�>� ��>�'�������F��G�����u�u�u�u�6�-����Y����VǶN��X���u��y�a�w�2����6����_	��
]�����6��'�2�`�[ϵ�	����K�N��D���4�%�0�9�w�$����T���F�=��Y��u�:�3�u��8�������X(��z��%���0�h�y�>�'�`�}��Y���S��V�����u�,�9�&�z�}�W���Aӵ��F��������0�6�:�<�o�W�������c��R	��Yʾ�%�h�_�x�w�}�W��*����V%�������x�_�x�u�$�<����Y����@"��V8�����u�=� �1�4�0�W������� ��ZN��ʺ�u�=�u����W��Y�ƨ�R��ZB�����u�=�,�4�2�3�Ϭ�T����@��R
��ʡ�0��8�9��6������ƴl�N�����!�4�u�=�w�8����
ӎ��VF��Z�����&�<�u�9�4�}����Y������CN��ʷ�0�_�x�u�#�.����ӑ��GF�������1�!�u�:�<�}�#�������R��R��ʼ�u�=�:�0�>�<��ԑT����Z��R
��ʡ�0�;�8�0�w�;�3���Aԕ��]F��T�����;�!�0�%�%�4����Y������Y	חX��� �0�{��6�9���Y����]F��U����� �%�'�9�:�)�W��s���2�������0� �%�!�1�4�����ƨ�A��[�����6�0�u�:�#�8����Ӄ��Q
����X���u�=�u� �'�)�Y�������R��RN�����:�%�:�0�#�)�ϒ�Y������P��U���8�!�<�_�z�}��������F��C����u�=�u����W�������Z��X��ʺ�!�:�u�0�2�s�W��s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߠ9�7�4�,�>�8�L�������V��D�����6�d�c�{�;�f�Wϫ�ӏ��VH��Z�����1�4�9�_�;�?��������9F��D������2�$�4�;�W�W���Y����6��s�����_�0�!�!�w�,��������V��Dd�����6�_�u��2�
����Y���\��YN�����'�'�;�0�f�}���Y���]ǻ�����1�=�u�u�w�g��������AF��Y	��D���:�d�u�h�f�f�Wϵ�����d��_N��U��<�u�;�0�2�}����Y����\F��T��F��u�>� ��4�����Y����Z��Y�����4�2�u�u�8�k�W��Y����F��G��U���u�u�u�u�w�3��������R��_����u�o�u�n�w�6��������F�N����;�0�0�u�6�:�W������\�N����!�_�u�4�'�8����Y���\��YN�����2�6�_�u�6�-����7���F������9�2�6�_�w���������F��T��ʦ�1�9�2�6�]�}��������F�N��Oʼ�u�!�
�:�>�f�Wϭ�����F�N��U��<�u�!�
�8�4�L���
����w��N��U���o�<�u�!��2����������R�����d�1�"�!�w�t�}���
����z��N��U���o�<�u�!��2����������C�����d�1�"�!�w�t�}���=����]W�N��U���u�;�&�1�;�:��������X"��V9�����u�:�;�:�g�f�Wϭ�����F�N��U��<�u�!�
�8�4�(�������w��`����1�"�!�u�~�W�W�������F�N��U���;�&�1�9�0�>�����Χ�R��^
��X���:�;�:�e�l�}��������F�N��Oʼ�u�!�
�:�>�����ۍ��G��S��Dʱ�"�!�u�|�]�}�3���0���F�N��U���&�1�9�2�4�+����Q����R1��C��U���;�:�e�n�w�.�������F�N����!�
�:�<��8��������d��_C����!�u�|�_�w�����N���F�T��ʦ�1�9�2�6�!�>����=����Z��_�����:�e�n�u�$�<����Y���F�N��U���
�:�<�
�2�)�ǵ�����W��N�����u�|�_�u��)�>��Y���F������9�2�6�#�4�2�_�������G�
�����e�n�u�&�6�<���Y���F��^ �����:�<�
�0�#�/��������[K��S�����|�_�u��#��F���Y���\��YN�����2�6�#�6�8�u�3���.����W��X����n�u�&�4�6�3�E���Y���	F����*���<�
�0�!�%�6��������F��@ ��U���_�u��!��l�W���Y�����D�����6�#�6�:�����������Y��E��u�&�4�4�9�i�W���Y����Z��C
�����
�0�!�'�<�<��������W	��C��\�ߊu��!��f�}�W���Y����]F��S1�����#�6�:�}��)� �������\��XN�N���&�4�4�4�>��W���Y�ƥ���h����_�u��!��)�W���Y���	����*���<�
�0�!�%�6��������[K��S�����|�_�u��#�����Y���\��B�����:�<�
�0�#�/����	����W��N�����u�|�_�u��)�8���Y���F���U���
�:�<�
�2�)�ǵ�����d��_C����!�u�|�_�w��������F�T�� ���!�
�:�<��8��������F��S��Dʱ�"�!�u�|�]�}�3���6����F�N��U���u�!�
�:�>�����ۍ��G��`����1�"�!�u�~�W�W�������F�N��U��� �u�!�
�8�4�(�������|��B�����d�1�"�!�w�t�}���=����F��N��U���u� �u�!��2����������C��"���=�d�1�"�#�}�^�ԜY����R)�� N��U���u�u� �u�#�����&����\��x�� ���1�=�d�1� �)�W���s�ƿ�R��B�U���u�u�u� �w�)�(�������P��������1�=�d�3�*����P���@"��V!��L���u�u�u�u�"�}��������E��X��:��� ��1�=�f�9� ���Y����F��V�� ��u�u�u�u�w�(�W���&����P9��T��]���!� ��1�?�l��������l�D*�����d�u�u�u�w�}��������T��A������!� ��3�5�FϺ�����O��N����� �d�u�u�w�}�W���Y����_	��T1�����}��!� � �9�������\F��d�����4� �d�u�w�}�W����ƿ�W9��P�����:�}��!�"�
����Hӂ��]��G�Uʦ�4�4� �d�w�}�W���Y����@��[�����6�:�}��#�(� �������\��XN�N���&�4�4� �f�}�W���Y�ƣ�GF��S1�����#�6�:�}��)���������Y��E��u�&�4�4�6�4�8���Y����\��D�����6�|�_�;�w�,��������V��=d�����0�!�'�u��}�ϛ�*����V ��C���ߠu�x�#�:�<�.�������K��X�����;�_�u�6�9�)����=����C��Y��U���;�0�0�u�j�i�W��MӠ��	��S��U���=�<�u�$�$�i�Y���s�Ư�]��Y��1���,�<�&��4�g�������F��A�����u�u�n�u�4�3����Y����G)��V��U���u�;�0�0�w�`����4����V��PD�����u�n�u�6�9�)����-����w��NN��U���;�0�0�u�j�6����	����VF�\*�����'�!�4�u�w�����4����9F��X �����>�8� �!�8�8����Y����T��S�����'�9�6�u�w�6����=�����������:�>�|�8�3�6��������9l�C�����4�u�,�0�8�}����Y����JF����ʴ�9�d�u�9�:�3�����ƣ�_��s��"���=�u�!�%�w�}����=����A��h��Uʼ�u�'�4�u�f�}�������\ ��C
�����
�0�!�'�<�<��������W	��C��\�ߠu�x�u��#��X���Y����G	��RN�����&�/�u�c�2�8����UӒ��Q��U�����'�%�'�,�%�.����Y���G��^ ��ʱ�!�{�u�3�2�}�����ƫ�G��E�����0�u�:�4�w�/����Ӎ��PF��MךU���;�9�&�4�6�3����Y���F�'�� ���!��'�,�#�g�WǱ�����N��_��H��r�|�_�u�$�:����=����]F�N��U���u�o��6�6�<�ǵ�	����W	��C��\���h�}�!�0�$�c�������A�dךU���;�9�&��#���������WF�=��1���
�}��6�f�9� ���Y���	[�X����}�!�0�&�i�m�^��Yӕ��]��D�����6�;��8�;�9�Mύ�����l��d��Dʱ�"�!�u�|�w�`�_������	��R��K��|�n�u�&�0�<�W�������_��V�����o�&�1�9�0�>�����Χ�C�
�����e�u�h�}�#�8����I����F��P ��U���0�=�<�u�w�}�W���Y�ƿ�W9��P��U���u�u�u�u�w�}�W��Y���9l�C�����'�u�:�u�.�>��������F��G��U���%�:�;�
�w�}�W���Y����A��F�����u�:�;�:�g�}�ϫ�
����WN��P\����>�#�'�9�4�t��������l�D�����&�:�;��4�>�W���Y����g��t�����o�u�:�=�%�`�_������V�UװUʦ�2�4�u�&�8�3�!���Y���F�N�� ���0�
�}��4�l��������\������k�:�=�'�j�z�P���s�ƿ�T��������6�9�e�w�}�W�������V������1�"�!�u�~�g�WǱ�����N��_��H��r�|�_�u�>�3�ϭ�:����e��[�U���u�u�:�;��>�ǵ�	����W	��C��\��u�:�=�'�j�u����
���O�=N�����9�&�� �#�8�3���Y���\��X��#���!�>�%�x�w�2����I����N��_��H���!�0�&�k�g�t�L�ԜY����R
��s��#���1� ��9�w�}�W���&����P9��T��]���6�d�1�"�#�}�^��Yۉ��V��	I�\�ߠu�x�u�%�4�<�W���Ӊ��\��B�����u�:�>�0�w�1�W������]����U���,�>� �%�#�4��ԜY����F��B�����4�'�4�
�w�}����������R	��U���2�u�k�u�1�.��������V��EF�� ���!�<�!�x�w�2����I��ƹ��Y�����4� ��9�w�}�W���Cө��C��V�����
�}��6�f�9� ���Y���F��C����:�=�'�h�p�z�^�ԜY����R
��s��:���u�u�u�u�w�}�W���	����G��E����u�:�;�:�g�}�J�������X��C����e�|�n�_�5�:��ԜY����V��G��1����u�'�8�>�9�����ƿ�T��DN�����'�4�u�3�$�+�Wϒ�Y����9F�N�����0�u�=�u�a�4��������@��V��U���u�!�&�8�4�}����Ӓ��D	��=N��Xʢ�!�u�=�u��<�����Ƹ�VF��D��ʡ�0�6�1�{�w�.�������F������e�_�u��#��;���P���@"��V'��N���&�4�4�;�0�o�W��
����z��=N��1�����}�|�k�}�3���0����F��V�����a�u�h�&�6�<���Yӕ��G��{	��\��u��!��b�W�W�������TN��R�����4�;�n�u�$�<�������[��s��<��_�u��!���_���E�ƿ�R��YV�Uʦ�4�4�;�2�n�}�Jϭ�����
]ǻ������}�e�u�j�.��������F��V�����d�|�i�u��)�>��B����w��~ ��]��u�h�&�4�6�3�E�ԜY����R/��PF�\��u��!��f�f�Wϭ������G��Hʦ�4�4�;�a�]�}�3���0����S�S��1����d�n�_�w�8����=����]\ǻ�����}��!���t�Wϼ���ƹF��X��U���e�!�u��4�l����s���F��V���u�h�}�!�2�.�I��P���F�D*������}��!� �9�������\F��R�����4�;�2������������Y��E��u�u�0�1�;�2�L�������A	��D�����%��!��l�W�W��Y����VF��RN�����,�6�� �#�/�[ϱ�Ӏ����_N��ǳ�9�0�{�u�?�.����
Ӓ��9F�N�����u�:�;�:�w�.����s�Ƌ�]5��T-�����&�_�u�:�w�}����Ƨ�C�	�����0�_�u�u�2��������F�������:�>�h�u�2�8����Y���K��_��*���#�'�9�6�>�:��������Al�N��Xǣ�:�>�4�>�!�/����?����AF��A�����_�u�u�u�z�5����Y����]��O(�����w�w�u�u�w�p��������a��CN�����u�u�u�x�!�2����;����_��V�����_�u�u�u�z�5����Y����A��E��U���u�x�#�:�<�<�8�������R��R-��;�ߊu�u�u�x�?�2�(���:������X��#���6�}�|�u�w�}�Z¨�����	��B �����u�%�;�u�w�}�Z¨�����	��D�����0�0�!�:�2�W�W���Y����P
��\��&���� �!�'�m�8����Y����)��E�����2�,�6�:�9�8�Wǌ�5���F�N�����6�8�%�}�w�}�W���YӍ��V��X�����'�h�u��2�>����Y���Z�^ �����o�u�_�u�w�}�W���:����~��V �����k�w�w�u�w�}�W���Tӏ����^ ��O���f�w�u�u�w�}����Y����l�N��U���4�0�0�u�w�}�W���Y����R
��N��U���u�u�u�x�w�3�W�������F�N��Uʗ�&��>�u�w�}�W���Gӵ��C
��[�U���u�u�x�u�9�}��������F�N��Uʷ�!�'�u�u�w�}�W���GӒ��VJ�N��U���u�u�x�u�9�}����������Rd��U���u�u��0��6�W���Y���X��V������y�u�u�w�p�W���Y����_	��Td��U���u�u�:�:�9�}�W���Y���X��D-�����6�6�}�|�w�p�W���Y����T����G���&�}��0�4�2�������F�N��6���!�4�<�u�w�}�J���	���F�N��U���u�x�:�!�5�2����Y���F������>�1�0�0�#�`�W������F�N��U���x�:�!�7�8�8����YӃ����R��ʒ�;�:�;�0�l�W�W���Y����A��dךU����0��0�4�2����*����\���� ���=�&�4�#�%�<��������T��EN�Yʴ�1�4�9�u�z�}�Ϫ�ӣ��P	�������u�u�<�!�w�;�E���<����@��_��U���1�u�&�%�3�4�Y���+����Z��X���ߊu�'�6�&��.����/����_Oǻ���ߊu�u�&�:�9�����H���	��R��Kº�=�'�h�r�p�t�}���Y����zF��^��ʾ�%�x�u�:�'�}�W���
����]��T*��D�}�:�g�0�$�u�8�������F��@ ��U���i�u�&�:�9�����Q����\��R��]���0�6�:�>�w�2����I��ƹF��Y
�����_�u�;�u�%�>��������T��B ��N�ߊu�x��9�.�)�ύ�����]����E���y�:�u�y�$�}��������R��T����� �u�!�!�2�}�Z����ƣ��������9�;�&� �w�8�����ƻ�G��=�����9�u�1�0�6�9� �������F� ��ʴ�&�;�=�:�8�.����Ӏ����Y�����2�7�6�u�8�)�ύ�����_��X���ߊu�9�� �#�8�M���	����@��V������|�u�7�0�3�W����ƾ�@��h���8�9��>�/�}����Y�����X��#���9�g�i�u�$�2��������l�N������0�6�:�<�n����s���F�D�� ���0��,�u�j�.�4�������_��=N��U���9�0�u�u�w�}��������P"��N�U���:�;��6�;�l�}���Y�Ʃ�WF��d��Uʰ�1�<�n�u�2�9��������_��B ����_�u�x��9�8��������|��T��ʼ�u�y�!�0�w�5�W���Y����]��XN�����"�9�u�0�e�}��������PF�������6�9�g� �8�W�������\"��V��U���9�0�u�u�w�}�W���Y����@%��Y�����d�"�0�u��2����=����[������u�u�u�u�w�}�Wϭ�:����e��[��ߊu�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}���Tӯ��F��V�����u�x�_�u�z������ƭ�C��E��ʼ�%�!�&�8�;�3�W����Ʈ�@��X ��:���6�:�>�u�w�/�D�ԜY����]F��S�����0�%�!�0�4�2�Ͻ�����TF��X�����0�9�u�:��0��������@l�C�����4�u�&�%�$�4���0ӑ��G��R�����#�'�<�;�w�;����������G��ʶ�1�{�u�x�w�8����Ӓ����E�����u�;�{�u�#�4�W�������\��U�����0�2�u�=�$�}����Y���G	��C��Yʷ�!�!�4�u�$�1����
Ӈ��F��RN�����&�{�u�_�w�8�>�������_�������3�>�#�'�;�>�J�������GǻN��X���:�
�u�$�9�(�$�������\ǻN����� ��8�9�9�o�������JF��E����� ��8�9�9�o����-��ƹF�	�����u�4�u�_�w�}�W���=����Z��S����4�<�!�y�w�p��������V��V ��U��!�u�m�o�w�e�W���Y����`��N��U��u��6�u�w�}�W��Y���Z��P�����0�d�!�u�a�g�W�ԜY���C	����U�ߊu�u�u�u�6�-����7���F�N��U���%�0�9��{�}�W���Y�������*���<�_�u�u�w�}��������F�N��U��u�&�:�;��>�W���Y���F���U���;��6�!�w�}�W���
����e��S'��U���u�u�k�&�6�<����0���F�N��Xʼ�u�&�1�9�0�>�W���Y����w��~ ��U���u�u�u�u�i�.�������F�N��U���x�<�u��4�<��������F��@ ��U���u�u�u�u�$���������^��SN��Kʦ��!��'�#�<����U���F��CN�����4�!�>�%�z�}�������	[ǻN��U���&�4�4�0�8�9���������V�����1�4�%�0�{�}�Zϱ�ӵ��w��h��&���d�1�"�!�w�t�M�ԜY���F��s��#���1�4�%�0�w�`�W�������_��V�����u�x�u� �w�)�(�������P������1�"�!�u�w�}�Wϭ�.����Z�N��U���u�k�&���<���Y���F�C����&�1�9�2�4�g�W��s�Ʃ�WF��Y�����0��%�!�6�-������ƓF��Y'�� ���8�9�;�f�4�W�W�������P
��\S����'�!�_�u�w�p����&�Ɖ�z��C=�����2�:�_�u�w�,����*����Z��X��U���<�,�"�'�y�,����*����Z��X��'���_�u�u�u�2�8�������F�N�����4�<�!�u�i�6��������F���U���0�0�u�4�0�}�OϪ�Y���F��=N��U���u��6�u�w�}�J���*���F�N��Xʼ�u�<�!�2�%�/����HӒ��P�
N�U���u�%�'�u�6�}�}���Y���`��[�����u�u�u�u�j�}��������KJ�N��U���x�u�;�u�#�����s���F�D�� ���0�u�u�u�w�}�J���
����G0��N��U���u�u�x�u�9�}����/����9F�N��U���!��9�1�9�}�W���Y����w��a�����u�u�u�u�w�p����
����\��=N��U���u��!��w�}�W���Y���X��s��<���u�u�u�u�w�}�W������C��C��]���6�d�1�"�#�}�^���Y�����V������8�9�1�w�c��������@��Z�����u�x�:�!��>����ۍ��PK��S�����|�o�_�u�w�}�W�������P	��d�����h�u�&�4�6�8��������WJ�C�� ���%��!�
���������\F��T�U���u�u�&��#���������WF�	N��1����9�1�4�'�8�[���T�ƣ�GF��S1�����#�6�:�}��>�FϺ���ƹF�N�����=�<�u�u�w�}�W���Gӕ��V%��^ �U���u�u�u�u�z�2�ϭ�����Z�
N��R���0�1�2�;�%�)�W���0����`��[��F���_�u�x�u�9�}����Y����_��=N��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�C�� ���<�!�'�y�8�8��������\ ��_��&���:�!� �&�]�}��������F��=N����� �%�!� �w�3�GϪ�Y����W��R �����_�u�u�x�?�2�(�������Z
��Ed��U���#�:�>�4�<�3��������}��N��Xǣ�:�>�4�&��9�4�������G��X	��*���!�'�&��"�)��������}��d��U���#�:�>�4�$�����?������V������8�9�1�w�}�Z¨�������V�����:�1�&��#�����*����VǻN��X���:�
�u��#��ϭ�����G*��!����� �|�u�u�z�+����ӕ��G��[�� ����!��9�3�(�;���6����G(��d��U���#�:�>�4�$�����������V������8�9�1��)�������F�A�����&���4�9�3����:����9F�+�� ���9�0�-�u�9�4�ϩ��ȉ�`��^������|�u�u�w�:����Ӌ��NǻN��U����0��1�?�}�W��Y����U1��C�U���u�x�<�u�>�)����C����9F�N��U���!��1�=�w�}�J���=����Z��N��U���x�<�u�<�#�:���Y��ƹF�N��:��� ��1�=�w�`�W�������Z��N��U���<�u�<�!�0�/�M���H���F������&�0��2�j�}�9�������A5��N��Xʼ�u�<�!�2�%�g�W��Y���F��d��U���u�u�u�h�w�����Y���F�C����<�!�2�'�m�}�}���Y���X)��E�����u�u�k�>�!�/����U���F���U���0�0�u�4�0�}�W���J��� l�N��Uʾ�;�0�u�u�w�}�W���6����G(��N��U���x�u�;�u�9�8����D��ƹF���ʸ�%�}�u�u�w�}�$�������F�N��H���4�%�0�9�{�}�W���Y���F�N��U���u�u�u�u�z�}��������T��N��U����8�9��<�%�W���Y����R��R-��;���u�u�u�u�w�}�W���Y���F�N��X���;�u�!�
�8�4�}���Y���@"��V��:��� ��u�k�$�4����6����G ��N��U���u�u�u�u�w�}�W���Y����]F��C
�����_�u�u�u�w��������F�S����3�:�1�u�w�}�W���Y���F�N��U���u�u�u�x�>�}��������9F�N��U���0��u�u�w�}�W��Y����U1��N��U���u�u�u�u�w�}�W���Y���F�C����&�1�9�2�4�}�W���Yӕ��V ��YN��U���u�h�u��2�����Y���F�N��U���u�u�u�u�w�}�W��Y���@��[�����_�u�u�u�w�.��������F�S�����4�;�u�w�}�W���Y���F�N��U���u�u�u�x�>�}��������9F�N��U���1�'�=�<��}�W��Y����_	��T1�����}�&�:�;��>�8�������O�C����&�1�9�2�4�+�}���Y���@��C�����;�u�u�k�$���������^��SF������8�y�u�w�}�W���Y����]F��C
�����_�u�u�u�w�.��������GF�S����!��'�!�6�-���Y���F�N��U���u�u�u�x�>�}�$���������N��U���&��!���>����Y����@"��V=�����4�%�0�y�w�}�W���Y���F�N��X���;�u�%��#��_���Y���F��s��:���u�u�u�u�j�}�3���6����_N��C��;���y�u�u�u�w�}�W���Y���F��CN�����2�6�#�_�w�}�W���=����R
��x��U���k�&�4�4�6�4�8����΃�G��y��\���u�u�u�u�w�}�Zϱ�ӕ��l
��^װUʰ�1�2�;�'�#�}��������F��=d��X���;�u� �u�>�)��ԜY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x�u�0�=�'�}�����Ƹ���DN�����:��u���W�W�������Z��CN�U���!��9�1�"����B���@"��V!��]���6�d�1�"�#�}�^��Y����R)��{������!��!�f�}����Ӎ��PO�
N�����&�k�:�=�%�`�P���P��ƹ��C�����h�&�4�4�"�u�^ǵ�����d��_C����!�u�|�_�w����������C����}��!� � �9�������\F��d�����4� �g�i�w��������X)��G�����x�u�:�;�8�m�L���
����|��R�����4� �}�|�<�(��������F��@ ��U���_�u��!��)�W��
����|��G��:��� ��1�=�f�9� ���Y����F��V�� ���i�u��!��)�B���6����G1��C��U���;�:�e�n�w�.�������F��V�� ���|�>� �%�#�4���Y����G	�UךU���!��!�u�j�.����������C��"���=�d�1�"�#�}�^�ԜY����R)��N�U���!��!�m������.����W��X����n�u�&�4�6�(�N��Y����R)��W�����%�!�<�!�z�}�������9F��s��:���e�i�u��#����Pۍ��G��`����1�"�!�u�~�W�W�������W�
N����� �}�d�}��)���������Y��E��u�&�4�4�"�l�W��
����|��\�����%�!�<�!�z�}�������9F��s��:���f�i�u��#����Pۍ��G��`����1�"�!�u�~�W�W�������R�
N����� �}�a�}��)���������Y��E��u�&�4�4�"�l�W��
����|��[�����%�!�<�!�z�}�������9l��Y
��!��