-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B+��t��ģ�1�x�u� �?�/�W���Y����Al�!�����9��:�0�#�}�/���L����9K�s��O���;�4�,�e�l�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����}�|�g�d�w�2�����Ƃ�G��V����� �0�!�u�8�-�������'��<������&�'�0�]�p�9�������z��E������!�'�4�w�3��������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��/����Y������G�����!�<�2�u�8�8����ӈ��Q��X������r�u�&�'�/�W���T���R��~<�����'�u��0�2�<�ϵ�����@6��d�����4�=�&�2�2�)�W���Y����9K�N�����!�u�;�!�2�>����YӲ��@F��C��ʺ�u��8�4�$�8�$�������~'��N�����u�u��8�6�.����ٍ��PL��A�����u� �7�'�8�}��������G�CחX����0�&�'�4�(�ϸ�Ӓ��@F��[��U���w�0�<�%�%�1����Y����Z��R�����9�'�!�u�z�}�W������T��YN��ʍ�9�;�u�<�#�%�CϚ�)ӓ��AF��^
��]���b�{�1�u�9�-�������KǶN��!���:�!� �u�$�.�4��� ����P	��DN�����=�u�� �w�;��������w5��+����6�;�x�u�w�3�ϼ�Y����V��GN��U���u���:�w�3����Y����#�CחX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�W�����ƥ�V��N��ʼ�0�{�!�
�8�4�(��M݇��l�B�����{� �0�<��)�Y���B���Q��NN����u� �0�"�%�s����W����9l������<�u�'�;�;�)�(���s����R��o�����'��7�_�>�/����7����l��RN��<���{�6�8�:�2�)�Y���B���@��_��ʡ�4�&�4�0�8�W�}�������B+��t��ʼ�u�_�0�0�>�u�Wϵ�����W��N��U��<�u�;�0�2�}�J��B���X"��V9�����u�u�u�u�9�4�������^��N�� ���6��'�0�w�}�W�������V�
N�N���>�%�u�u�w�}�W���Y�ƥ���R	��U��d�_�u��2�>����Y���\��YN�����'�'�;�0�e�)�W���D���l��E��Uʆ�8�9��>�w�}�W���Y����G��X	��N����8�9��<�%�W���Y�ƥ���h����_�u��0��<�W���Y�����D�����6�_�u��2�
�W���Y���\��YN�����2�6�_�u��8�3���Y���F������9�2�6�#�4�2�_�������G�
�����e�n�_�u�$�8����0���F������9�2�6�_�w�.��������]F�T��ʦ�1�9�2�6�!�>����Y����G	�UװUʦ��!��9�3�3�W���Y����G��X	��N���&��!��w�}�W���Y�ƥ�5��s��*����6�d�1� �)�W���s�ƿ�w��V��:���u�u�u� �w�)�(�������P��Z����!�u�|�o�w�2����D����]ǻ������9�1�u�w�g����
����\��d�����6�8�9�!�w�}�W����ƿ�W9��P��O���e�u�n�0�3��:�������9l��E����� �0���8�}����:������=N��X���:�
�<�&�6�)�W������l��R �����:�&�4�!�<�(�:���Y���F�T�����0�u�h�>�"���������X5��dךU����0���w�3�ϰ��Ƹ���R�����0�4�u�3�<�(�:���T�ơ�P�D��ʡ�0�0�u�x�w�.�P���Y����Z��V�����"�!�u�=�w�<�ϳ�����R��Z�����4�1�9�,�8�}�}�������]��z�����u�u�u�u�w�}��������N��B�����|�d�_�u�z�}����Y����5��Dd�����u�;��!��1�Ϸ�Y����JF��z�����x�u�:�;�8�m�W���
����\��h�����>�4�4�<�#�p�W������]ǻ��ʔ�9�4�4�'��}�Ͽ����X5��_�����:�d�u�3��8��������9F��^	��ʦ��9�4�4�%�.�W���Y����_
��C�����o�u�:�=�%�`�_������	��R��K��|�|�_�u�#�-�W���=����R
��d��ʼ�u�'�4�u�<�<�3��� ����\��XN�U���&�1�9�2�4�W�W���ӧ��w��a�����
�u�&�4�%�$�_�������\��XN�U����0�4�4�6�4�$������@��V������!��9�3�/����Y����R��V��&���!�o�u�:�?�/�J�������X�G����x�u�<�;�;�}��������]��R�����=�u��&�w�)��������R��CN��U���4�u�>� ��>�W������F����*���<�
�0�!�%�6��������F��@ ��U���_�u�<�;�;�.�3���:����z�N��U���4�4�=�<��}�J�������X��C����e�|�n�u�$�:����
����p��Y!��U���u�o��!��<����C����G��DS����'�h�r�r�~�W�WϪ�	�ƍ�W��V��ʼ�u�'�4�u�<�(�:���Y����G	�N��U���
�:�<�
�2�)�������\F��d�����4�u�&�1�%�5����Y���F��v
��6���;�!�o�u�8�5���Q����A�^��\�ߠu�!�%�u�4�(�4�������@F��E��]���8�4�&�1� �)�W����ƿ�W9��P�����:�}�b�1� �)�W���s�ƿ�T��������4�;�u�w�}�W�������[��h��H���!�0�&�k�8�5���^���lǻ�����&��!��;�9����0�����h�����0�!�'�>�"���������V�S�����'�h�r�r�l�}�����ƿ�w��a�����<��!�o�$�9��������G	��\ ��8���u�:�;�:�g�}�J�������X�G�Uʦ�2�4�u�&�2�5����Y���F�N�����2�6�#�6�8�u�9�������\��XN�U��}�!�0�&�i�m�^�ԜY����R
��D/�� ���9�1� �u�w�}�W���&����P9��T��]���8�4�&�1� �)�W���C����G��DS�E���_�u�<�;�;�.� �������JF�N��U���!�
�:�<�w�`�P���s����Z��[N��6�����'�,�w�}�W��
����\��h�����>� ��6�z�}�������	[�X����r�r�n�u�$�:����
����r��N��U���u�o�&�1�;�:��������F��@ ��U���u�u�u�u�w�`�_������V�d�����4�u�&�:�1�<����Y���F��D�����6�#�6�:��j��������F�N��U��}�!�0�&�i�m�^�ԜY����R
��D"������0�&�u�w�}�W���&����P9��T��]���8�4�&�d�3�*����P���	��R��K��|�_�u�&�0�<�W�������_��{��U���o�&�1�9�0�>�M���I��Ɠ9��^ װU���u�=�u�:�1�����Y����@F����U���2�4�8�;�w�4����Y����*��q>��Yʴ�1�6�0�!�$�}�Z�������@F��EN��ʐ��6�-�6�:�2�����Ƽ�\��ZN��ʶ�0�3�6�0�#�4�������K��^�����0�u�4�_�w�p��������B%��Q"�����u���0��<����Y����G��X��0���0��4�0�w��;�ԜY�ƫ�]��TN�����u�u�u�>�!�/����Y����|��T�����x�u�;�u�9�8����D��ƹF������1�=�h�u��8� ������F��N�����'�o�u�m�w�}�Wϵ�����@F�
P��;���4�&�u�u�z�}��������AF��_�U���%�'�u�4�w�W�W���Y����_��\N��U���k��8�9��6�W���Y�������*���<�_�u�u�w�<��������F�	N������>�-�u�w�}�ZϷ�Yӕ��l
��^ךU���u��0��6�}�W���D�ƿ�\��X��U���u�u�x�<�w�.������ƹF������u�u�u�u�j�}�4���.���F�N��Xʼ�u�&�1�9�0�>�W���Yӕ��V ��YN��U���h�u��0��3�W���Y���F��N�����2�6�#�6�8�u�4���.����W��X����_�u�u�u�$�2�������[�D�����1�y�u�u�w�p����
����\��h�����d�1�"�!�w�t�W���Yӕ��\��R/�����h�u�&�:�1�8����U���F��CN�����2�6�#�6�8�u�9��������Y��E�ߊu�u�u�&�8�;����Y���F��t��1���y�u�u�u�z�2�ϭ�����Z��R��¾�:�3�<�!�z�}�������F�N��9���<�2�:�3�w�c��������p	��DG�X��� �u�!�
�8�4�(�������}��V��Dʱ�"�!�u�|�]�}�Z���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǻC�"���u��6�d�w�5�W���Y����]F�������<�!�u�0�:�3����<����@��R ����� �0�_�u�z�<����
����UF��RN�����6�0�!�{�w�5�W��������������0�u�:�0�?�/�W��Y����R
�������u�;�'�&�"�>�ϼ�Y����Z��PN��ʦ�<�!�<�u�9�8��������GHǻC�0���u�0�8�;�w�8�Ϸ�^�ƥ�C��S��U���8�4�1�3�2�8�Ϸ�	���@��RN�����4�0�u�x�w��Ϸ�	����F��_��U��� �&�=�#�w�2��������WF�������=�u�<�0�>�8���� ���F����U���#�:�&�&�0�8�������[��^����� �<�2�<�1�/����+���l�CךU���u�u�u�u�w�}�W���&����lF�N��*���
�u�u�u���(���Y���F�N��U���u�u�u�u�w�}����Y���F��N��	���u�u�u�u�w�p�W��������C��U���&�)�x�x�w�<�Ϣ�T�˰�~���X���{�u�x�u�w�}�W���Y�����h1��	���x�
�
�
�+�}�Z���&����F�N�U���u�u�u�u�w�}�W���&����N��U���u�_�u�x�w�}�W���Y���F��N��U���)�u�u�u�w�}����T���w��~ ��\���x�u��d�+�p�W���Y���F��N�U���u�u�u�u�w�}����&����F�N��U���u�_�u�x�w�}�W���Y���F��h1��*���u�u�u�u�w�}����T���F�N��U���u�u�u�u�+�}�W���Y���F��N�U���4�4�;�/�w�p�ύ�5�ư�K�C�X���x�u�x�u�w�}�W���Y�����h1��	���x�_�u�x��>�W�������E��e"��ʹ�;�0�y�!�w�<�����ƥ�P��D�����,�:�u�=�w�<��ԜY����]	��R�� ���u�=�;�u�$�)�Ϛ�����Z�*�����<�u�&�4�$�}�����ƥ���=N��Xʆ��u�9�;�w�4�Ϫ�ӂ��RJ��XN�����!�9�;�&�"�}��������[��^ �����u�;�:�u�z�}��������V��Y����x�u�x�u�6�5��������\��^ ������6��'�2�}����YӲ��A��E��&���&�2�0�!�y�W�W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��=d��X���=�&�u�'�6�.��������VF��C��'���u�&�1�!�w�8�����ƨ�G��X�����;�y�_�u�z�n��������V��Y��Uʆ�:�;�4�u��l����*����Z��U��U���2�4�{�u��1�M���	����@��V������|�u�7�0�3�W����ƾ�@��h���8�9��>�/�}����Y��� ��'����!�u��6�f�1��ԜY���F��EN�����u�:�>�4��1�������F�N��Uʼ�u�h�u�=�9�}�W���Y�����[�����9�}�|��w�`��������zO��s��"���=�d�1�"�#�}�^�ԜY���F�N��4���4�4�4�<��1�_���3�����V������n�u�u�w�}�Wϻ�
���F�N��Uʦ��9�4�4�%�.�>���P���@��[*�����&��}�x�~�6��������F��@ ��U���_�u�u�u�w�}�W�������R0��^
�����|��u�h�$���������W5��DF��]���|�_�u�u�w�}�W���Y����F�N�����9�:�n�u�w�}��������9F���U���_�u�;�u�%�>��������9l�C��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�u�x�w�5�Ͻ��ƭ�G��R�����4�4�u�4�6�<���.����]��S
�����=�u�4�u�2�0����Y���C��C�����<�2�4�:�2�}�Z�ԶYӕ��P��t����u�h�}�!�2�.�I��P���@��S�����e�u�i�u�$�9��������9F��D9�����}�|�u�u�j�.� �������lǻ/�����4�4�=�<�m�}��������@"��V-�����!�u�&�4�6�3�W�������R5��DB�����4�4�<��6�3���s���F�N��1����9�1�;�w�.��������Z��[��Uʷ�2�;�_�u�w�p�����ƣ�VF��P�����=�<�u�4�6�(�W�������W��^ ����u�u�3�'��4�W���Ӎ��^+��DC����_�u�u�u�$�<��������zM��R�����!��4�;�"�u�^�ԜY���@��C�����=�<��}�|�t�K���
����e��S-�����!��n�u�w�8�ϲ���ƓF�C�����4�;�e�u�$�5����Y����\F��RN�����&�2�0�!�w�}��������Z��^��I���&�4�4�;�g�u�3���.����W��X����n�u�u�&��)�!�������]/��G��Hʦ��!��9�3�3�}���Y���@��C��]���<�u�0�4�2�}����������C�����;�u�0�8�9�W�W���Tӕ��R��YF�U���1�9�,�1�6�9�����ƹ���C��F���&�2�0�!�w�)�}���Y����yF��_��ʾ�%�x�u�:�'�}�W���
����R%��^ ��]����8�4�&�2�����D���F�N��4���4�4�'�&��u�]�������c��R	��\¾�4�4�<�!�z�}�������9F�N�����4�4�<��6�3�ǔ�����R��R�����h�_�u�u�w�}����=����R
��d��]����>� ��4�����T����F�R �����n�u�0�1�'�2����8����["��V-����_�u�x�u�z�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��ƓF�-�����3�>� ��4�}�6�������F��Y#���ߊu�:�u�u�9�m����7����P�	�����0�_�u�u�z�5����Y����P(��N��Xǣ�:�>�4�>�>�.�>����΅�^	��\ ��8����'�0�|�g�}�W������l��q�����=�<�u�h�]�}�W�������RF��t��"���&�:�3�0�%�<�_���Y�����X��U���:�1�;��2�.��������p	��DF�����u�x�=�:��}��������@"��V-�����}�|�u�u�z�+����ӕ��R��B�����4�=�<��#��}���Y�˺�\	��VN��1����9�1�;�$���������R��YF�����u�x�=�:��}��������W)�������4�<��4�9�(�_���Y�����X��U���4�4�0�;�$�
�4���ۯ�F�C�����4�&��!� ��ϭ�.����Z��_��U���x�#�:�>�6�.�6���������S
�����}�|�u�u�z�+����ӕ��W��D��ʦ��1��4�9��F�ԜY���E��\1�����6�8�;�&��>�����΅�9F�C�����
�u�&�6�"��ϭ�8����p��YF��D�ߊu�u�x�=�8��W�������R
��x�����6�8�4�<��)�>�ԜY���E��\1�����0��!�:�2�W�W�������K��R �����:�>���4�%�_���P���F��R �����4�u�_�u�w�}�W�������p��YN��U��y�u�u�u�w�}�W���Y���F�N��Uʷ�:�0�;�o�w�<��ԜY���F��^��<���2�u�h�u��0�ϵ�����@6��d��H���u�x�<�u�5�2����C�ƪ�_��N��U���>�:�3�<�#�}�W��Y����U1��C�U���u�u�u�u�w�}�ZϷ�Yӏ��V�������m�!�u�m�m�}�O���Y�����C�����u�u�k�>�6�<����U���F�N��U���x�u�;�u�9�8��������^��XN�U��d�_�u�u�w�}�8�������F�
P��:���6�:�>�u�w�}�W���Y���K�^ �����2�'�'�;�2�o����Y���9F�N�����8�%�}�u�w�}�Wύ�����_��N��U���8�9��<�%�W���Y���F�C�����!�
�:�<�]�}�W���Y����V ��S��U���h�u�&�:�1�9����Y���F�N��Xʼ�u�&�1�9�0�>��������W	��C��\���u�u�u�&��8� ���Y���[�D������'�,��{�}�W���Y����]F��C
�����_�u�u�u�w�.�������F�
P�����3�4�4�u�w�}�W���Y���F��N�����2�6�#�6�8�u�4���.����W�N��U���&��4�<�0�2����D�ƿ�	��^ �����}�|�u�u�w�}�ZϷ�Yӕ��l
��^ךU���u�u�&�4�6�3�W���Y�����V������}�|�u�w�}�W��Y���@��[�����6�:�}��#�
����H���F�N��1����!�u�u�w�`�W�������R��B��\���u�u�u�x�8�)��������l��C�����4�<�!�x�w�}�W���Yӕ��R��V��<���u�k�&��#���������]N��N��X���;�u�!�
�8�4�}���Y���@��C����� �u�h�u�$�<��������Z��CF��Y���x�:�!�&�3�1����Y���F��D*�����;�u�u�u�i�.� �������J�N��U���u�x�u�;�w�)�(������F�N��1�����!�u�w�`�W�������]N��G�U���u�u�u�x��)��������9F�N��U���1�'�&��w�}�W���
����A%��^ ��\���u�u�u�u�z�}��������T��A�����u�:�;�:�g�W�W���Y�ƿ�r��R�� ���u�h�u�&�3�/����Q����F�N��U���:�!�&�1�;�:��������F��@ ��U���o�u�u�u�w�.�6������F�S����6�8�=�<��t�W���Y���K��YN�����:�<�
�0�#�/�C�������V�N��U���&��0��#�}�W���D�ƣ�V�N��U���u�u�u�u�w�}�Zϱ�ӕ��l
��^�����'�a�u�:�9�2�G�ԜY���F��v�����u�u�u�h�w�.����:����/�B��U���u�x�:�!�$�9��������G	��Y�����:�e�_�u�w�}�W�������R
��x��H���&�6� ��;�9����P���F�N��ʦ�1�9�2�6�]�}��������G��R ����_�u�&�&��/����Y����@'��B�����>� ��6�~�W�W�������R
��N�U���6� ��9�3�(�_�������W�=d��:��� ��o�u�'�2����*����V%��y��Uʷ�2�;�u�u�>�}��������VN��Z��6���-�u�=�;�w�}�Wϭ�.����Z��NN�U���0�=�<�}��0����B���F��D/�� ���4�0�6�u�j�3�ϭ�.����Z��NUךU���;�u�3�_�w�3�W�������|��B��N�ߊu�x�6�0�#�}����������CN�����!�0�4�6�:�1��������G	��T�� ���0�4�1�"�2�W�W���ƿ�R��X��[���=�u�0�4�w�.�������� �������:�>�u�u�$�}�}���
����^��C��Hʦ��6�8�9�#��ϩ��Ƨ�E��[��H���9�0�;�!�$�
�4�������9l��SN��9��