-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����9�6�{�=�]�p�6�������\��v�����y��&�u�2�)��ԑTө��T��[N�����!�u��0�b�i�%��Y����	F��$����d�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��ƴF��N�D���:�,�<�=�w�<����ӯ��G��R ��U���%�'�!�:�]�p�6���+����@F��D���߇x��!�:�6�}��������@F��C�����;�:�8�!�8�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��CחXʅ�'�:�0�u��4�W���Ӆ��R����ʺ�u�=�0�u�%�>����ӓ��G��X�����'�6�<�;�;�p�W���Y���F��T�����u�4�=�'� �2�W�������]��Y��U���4�%�:�0�$�3�W�����ƴl�N��U���u�u�&�u��0����������D�����=�u� �7�%�2�W�������]��Y�����u�:�7�_�z�}�W���Y����A��R
�0���u�'�6�&�>�:����	����A��T�� ���<�;�u�;�2�8����Y����9K�N��U���u�0�6�u�#�8�W����ƣ��������'�!�:�u�2�}�ϭ�����[��a������4�!�=�$�W�Z���Y���F��Y
��'����1�0�&�9�p�}��Y���F�+��ʥ�:�0�&�;�w�1����������R�����9�!�:�u�!�/�W���ӕ��R��_��#���1�x�u�u�w�}�W���
����@H��CN�����=�;�6�9�"�<�Ϫ�Ӏ��G��X�� ����6�8� ������Y��ƴF�N��U���#�9�1�"�2�}�6�������R
�������{�x�_�x�w�}�W���Yӳ����C��4���<�0�!�u�9�4��������Z��X������!����<�ϭ�����e��S@חX���u�u�u�u��*����Y����[��R
�����!�0��!�w�8�����Ƹ�VF��E��X���u�u�u�u�w�/��������]��^ �����7�:�>�7�w�.�����ƿ�R��Y8�����<�=�#�9�3�p�W���Y���F��C��ʦ�4�4�;�z�y�	�ϗ�	����R��^�����1�7�u�9�w�5�W�������]��[���߇x�u�u�u�w�}�$����ƿ�^�������4�0�&�%�8�)�ϼ�Y����A��PN�����;�u�9�8�9�}�Ϫ����F�N��Uʦ�4�4�;�4�>�}����s��ƴF�N��U����!�u�&�3�1����������*��ʗ�3�0�&�u�?�$���� Ӓ����R�����;� �u�4�6�p�W���Y���F����U���&�u�<�&�{�<�����ƨ�_��T�����!�&�3�'�#�8����Y����V��YN����� �_�x�u�w�}�W���	����@��PN�����u�0�:�1�w�}��������V
�������4�0�u�:�w�5�W���	����Z	��C��U���u�u�u�<�2�.�����Ƹ�VF��R�� ����{�x�_�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9
��E��U���0�u�:�>�]�}��������G��X	��*��a�4�9�_�w�.�W���݈��V��h��[���n�u� �0� �/�Y���?����Z	��[*�����:�{�9�n�w�(�ϩ��Ȝ�T(��C������%�4�9�]�}��������X��G@���ߊu�&�u�:�<���������p	��Q�����{�9�n�_�>�/����7����l�B�� ����{�6�8�8�8������ƓV��C������6�'�6�;�>�W���YӁ��V��d��Uʾ� ��:��8�6�W���ӏ��V��N�U��u�u�>�4�6�3��������Z��Y�����4�2�u�u�8�o�M���P���C	��d��Uʦ�&�'�0�0�w�g��������]]ǻN�����0�9�u�u�9�.��������9F�������0�3�o�>�}������ƹF��g�����'�8�;�u�w�3��������X(��g�����&�d�1�"�#�}�^���T޳��W��N�����6�,�9�&�>�(�8���Cӏ��F��P ��]���:�;�:�e�l�}�Z��A���F��C��%���0�4�<�u�w�3�5�������P�������6�9�6�&�z�l��������l�N������4�0�o�>�}����8������Z>�����6�&�x�d�3�*����P���3��_�U���&�0�1�1�%�.�>���Y����]��Y��4���!�>� ��8�����T�ƨ�D��^�U���l�l�_�u�w�p�6�������A	��D��ʷ�:�>�u�=�%�}��������R��=N��U���!���9�3�g��������]0��C�����4�;�'��-�}�W�������V�=N��U���!���o�>�}�����ލ�A��CF�����;�'��/�w�}�W������]�=�[�ߊu�u��!���MϷ�Y����V��v�����>�4�4�;�%�����Y�ƨ�D��^�U���d�{�_�u�w�p�W���Y����F��V�����&�0�0�u�9�}��������\��_�����u��6�8�"�����CӉ��$��[��#���:�}��8�%�>����
����\��XN�N���u�&�6� ��)�W����ƈ�G��C/��*����8�'�6�;�>�������\F��N��X��{�_�u�u��>����(����F��V�� ���,�!�>� ��2�5�������W	��C��\��u�x�a�{�]�3�W�������c��u���ߠ4�6�<�0�#�/�W���Y����A��s�����9�6�u�&�]�}����*����WR��E��U���4�'�,�u�6�(��������X������0�}�b�1� �)�W���s�Ƹ�C��Y�����g�'�
�u�$�<����Y����A��E����u�u�3� �$�:����Hӂ��]��G�Uʡ�%�u�;�<�9�9�6���ӏ��R��NF�����4�u�4�2�w�c�^ϱ�Y����T��Y�����:�e�n�u�#�-�W�������V��S/��*���&�4�'�,�w�<����Y����VF�G��ʀ�&�2�0�l�%��_�������q
��\��U���;�:�e�n�w�)��������W'��h��ʴ�'�,�u��:�/��������Z��S�����|�:�u�=�$���������A	��[����1�"�!�u�~�W�W���Ӥ��_��a������!�<�u�%�<�_�������V��Y	�����1�"�!�u�~�2�W�������V��EF�� ���:��:�>�z�}�������9F��N��7���0�;�0�!�%��(���
Ӈ��R��y�����&�<�2�;�#�}�W�������V�X�����4��6�:������8����I�
�����e�n�u�!�'�}����K����l��DN�����>� ��:�2�.��������\��XN�U����2�0�a��$�ǵ�����P$��T��Dʱ�"�!�u�|�]�}����*����WW��E��G���u�&�4�'�.�6��������Z��Y��U���;�:�e�u�1�����H˧��R��������,�<�0�f�9� ���Y����9F��^	��ʦ�4�4�4�<��$�MϜ�����e��X��7���o�u�:�=�%�}�I�������[�Q�����_�u�<�;�;�.�������5��Y��M���4�g�
�n�w�.����Y����R'��fN�&���0�d��'�.���ԜY����R
��g�����<��'�,�m���������\��v1�����<�;�9�&�?�.�6��� ����[��
�����_�u�<�;�;�.����/����r��NN�7���0�;�0�!�%��(��Yӕ��]��D/�� ���'�,�u�u�4�(�E��� ����F��P ��U���6�8�'�4��g�6�������J9��=N�����9�&�6� ��)����0����P��
�����_�u�<�;�;�.����6����A��T�����g��,�!�]�}����ӕ��R��S�����4�u�u�0�3�9����K����l��y�����&�<�2�;�#�}�������9l�D������"�&��2�;����?����Z��tN� ���2�0�d��.�)����)����@��P;�����u�u�:�;�8�m�L���
����_F��^	�����0�3�;�0��/����8����f��P ��Dؔ�,�!�>� ��2��������G�
�����e�n�u�&�0�<�W�������A��~ �����u�0�1�1�%�.�E��� �����Y��E���h�}�!�0�$�`�WǱ�����X�X�����k�r�r�|�l�}�����ƿ�@��C-�����%�u�u�:�;�<�!����Χ�F��X����� �<�&�1� �)�W���C����G��DN��U���&�|�_�u�4�3����Y����w��u�����o�<�!�2�%�g�W�������V��Y	�����x�d�_�u�>�3�ϭ�����U)��a�����:�9�4��4�2�_�������q��R��Dʱ�"�!�u�|�]�}����ӕ��G��Q!��<���<�;�1�m�%�o�(���7����G��Q����1�"�!�u�{�6��������Z��N�����u�|�_�u�>�3�ϭ�����U)��fT�����1�m�'�g��u�9�������U ��DC����!�u�y�>�6�<����*����F��@ ��U���_�u�<�;�;�.��������	F��D������9��6�2���������]��T��]���0�&�h�u�g�t�W��,����F��P ��U���%�9�;��;�$����<����	F��D������9��6�2���������]��T��]���0�&�h�u�g�t�}���
����_F��D������%�o�7�8�8���Y����l�D������&�!�0��4����Cӄ��_��T�����0�_�u�<�9�1��������c	��C��%���o�7�:�0�9�g�W���
��ƓF�A�����2�!�'�_�w�p����&����]ǑN�U���0�9��0�1�4�Ϻ�����^�������{� �0�4�<�8�W���Y�ơ�K9��Y��U���=�9�u�=�w�2��ԜY����V��C�����;�u�'�#�9�}��������^��^ �����'�9�7�:�<�}�������F��C�� ���>�0�u�u�#�4��ԜY����Z��RN�����3�&�&��#�2����	����Z��[N��Uȡ� �w�_�u�z���������[��q�����u�:�=�9�w�4�Ϫ�����R��Y�����0�{�u�4�#�4��������\ ��u�����/�u�u�<�9�1��������l�V�����0�>�0�u�1�.����4����Z��E����&�2�4�u�$�����B���R��^��ʸ�-�3�;� �m�.����B����G��U��U���
�4�:�!�8�}�"�������U ��G��Oʦ�2�4�u�&�u��}����ƓF�=�����!�0�6�'�2�)�;���
����U ��S�����<���4�3���������U/��R�����&��u�4�"�.�W��Y����WF�������4�0�3�9�2�}�Ͽ�ӓ��]�N�����&��8�9��6�}�������F�^�����2�0�2�}�6�-����PӒ��]l�N�U���<�u�8�:�#�3�W�������@3��v�����u�&� �0�w�3��������C
��R����=�"� �1�4�8����s���K��B	�����:�!�u� �w�8�����Ʃ�C��������0�3�!�w�5��������\ ��Y@��ʼ�u�=�;�0�]�}�W���ƻ�_
��RN�����0�u�,�&�!�/�Ͻ�����\ ��V�����,�'�&�!�>�:�W���
Ӂ��V��Dd��U���u� �1�0�$�2�W�������\F��X�����!�0�&�9�4�4�ϱ�Y���� ��C��6���3�6�0�!�w�.��ԜY���1��C��U���4�!�2�u�1�)����	����P��R��ʥ�%�9�;�u�?�}��������\F��S��U���u�4�x� �]�}�W���Ư�V��Y	��U���<�u�3��y�
�W���Y����JF��_��3���;�0�6�u�2�8�����Ƥ�_��_��4�ߊu�u�x�!�8�.��������W��V �����>�8�8�'�2�}�Ϫ��Ƣ�V��X@ךU��� �0�9��2�;����E�ƿ�@��C-�����%�}� �0�;���������Z��N�����u�|�s�&�$�������ƹF��Y
���ߊu�;�u�'�4�.�L�ԜY����V��X��<���-�:��<���G���DӒ��F��P ��]���"�&��0�1�3��������~��[�D���"�0�u� �2�1�4�������W�N��U���u�u�u�u�w�}�W���Y�����RN�����&�2�0�}��*��������W��X������y�g�n�]�}�;���
����U ��S�����<���d�w�`��������V��{�����0�3�;�0��/��������J��N����� �0�9��2�;����H���F�N��U���u�u�u�u�w�}�W���������B �����}��"�&��8��������g��z/��Y��n�_�u�� �.�4�������K ��c��8���g�u�h�!��3����ۍ��D��t�����0��'�=�$�<�6���U���D��������0�3�<�2�l�}���Y���F�N��U���u�u�u�u�w�8��������@��R
��9���&��0�3�9�8�1�������pT�G�����2�0�!�8�;�>�������[��v-��\��u�:� �&�0�8�_�������p	��Q'�����'�=�&�4��)�[��Y������R/��6���3�<�0�d�]�}�W���Y���F�N��U���u�u�u�0�$�}��������V�������:�3��1�/�2�#���4����T�=d�����=�&��0�1�3��������~'��G��Hʡ�
�;�<�;�3�6����
����U ��S�����<��6�9�f�l�^ϩ��ƿ�@��C-�����%�}�|�u�w�}�W���Y���F�N��U���u�u�9�0�w�2��������X.��_��6���3�;�0��%�5����H����lǻ�����!�:�3��3�%��������T�S�����&�2�0�}��:��������]��q�����4��!�y�e�}����
����_��R�����d�_�u�u�w�}�W���Y���F�N��U���0�&�u�!��3����ۍ��T��C-�����1�-�:��>��4��K��ƓF�>�����0�&�0�1�3�/����Y������T�����&�!�u�:�'�3��������[��_��U���9�u�0�!�%���ԜY����]��V������!�4�<�w�4����ӂ��R��C�� ���!�0�3�'�#�-����
����Q
��\d��X���'�6��6�%�>��������_F����ʴ�u�=�u�"�w�$��������]��R��U���!�0�0�&�0�<�ϼ�����F���ʴ�0�&�;�u�8�)�ϸ�����A��s�����0�:�,�7�8�6�}�������@N��Z��6���_�u�0�<�]�}�W�������T9��P�����0�9�|�!�2�W�W���Y����W'��E��<���%�u�h�&�2�9����
����Z��D<�����'�&���'�z����Hӂ��]��G��U���4��1�0�$�3�}���Y����Z ��N��ʥ�:�0�&�_�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�}�Z�������w��,�����o�u�x�u�?�/�W���Y����X��DN��U���4�!�4�u�?�}����Ӊ��G��SN�����&�;�u�;�#�}����T�Ƣ�GF��R
�� ���2�4�6�9�"�<��������[��V�����&�4�!�1�]�}�Z���Y����R��G�����;�u�;�!�6�)�Ϫ�Ӏ��@��Y�����&�!�0�6�;�(����Ӈ��F�N��U���u�4�4�:�1�8�W���Ӕ��C�������%�0�<� �w�/��������]��:��U���4�u�x�u�w�}�W���ӏ��G��Q��ʥ�:�0�&�;�w�3�Ϸ�Y����]��R
��ʡ�0�&�6�;�w�3�W������K�N��U���6�&�<�2�"�4�Ϸ�Y����P��R ����� �4�<�;�w�5�W���ӈ��W��U���ߊu�x�u�u�w�.����Y����V��Y	�����<�u�:�u�2�9�ϱ�Y����G��SN�����&�;�u�;�#�4�}���T���F��_�� ���;�u�4�6�;�)���Y���F�N��ʱ�!�u�3�&�#�?����Ӗ��P��^ �� ���&�<�u�$�6�}�ϭ�����P
��d��X���u�u�u�<�4�}�����Ƹ�VF��Z��U���&�8�9�&�"�8�W�������[��V�����:�u�;�u�z�}�W���Y����C��^��U���!�_�u�x�w�}�^ϊ�Ӣ��RF����U���:�1�4�1�#�4�ϫ�����@F��[�����1�:�6�u�?�W�W��Y�����A��ʥ�:�0�&�;�w�3�ϸ�����@F��DN�����3�!�0�6�;�(�������K�N��U���u�8� �!�8�}��������V
���� ���1�!�u�:�'�3��������[ǻC�U���u�6�8� �6�4�Ϫ��ƿ�V��^ ��U���#�:�&� �>�}�ϭ�����P
��d��X�ߊu�x��u�6�}����Y����G�������1�1�!�u�"�.����Ӓ����T����� �<�&�!�]�}�ZϺ�����VF��RN�����'�$�<�0�w�3��������^��E��[ʁ�0�1�!�u�$�.����s�����S��U���3�'�u�=�#�<�ϭ�����R��D�����=�u�'�6�"�4�W���
ӏ��G��=N��Xʰ�!�!�{��2�8�����ƨ�G��B��ʷ�!�0�;�&�6�<����Y����G��D���ߊu�x�%�:�2�.��������]�������7�3�0�u�2�*�����ƪ�A��U�����;�u�=�_�w�p����Ӗ��P��^ �� ���{�u�x�_�w�p�#�������^��E��U���u�!�'�u�f�}�&ϭ�����F��R �����'�6�;�!�w�p�W���������T�����u�!�6�;�"�8�W���(ӕ��C
��R��ʶ�6�0�_�u�z���������@����ʻ�0�&�&�4�4�$����
����V��XN��U���<�4�9�_�w�p�����Ƹ�VF��V�����&�:�u�:�'�)����Y������C��ʳ�'�0�6�_�w�p��������\�r��U���4�8�8�'�w�8����ӎ��WF��RN�����,�9�&�u�z�}�����ƥ���S�����!�0�1�!�w�)��������E��B��ʡ�0�&�4�6�.�1����T�ƥ���Y
�����=�u� �'�9�}��������]HǻC�1����8�'�u�2�(������� L��V��6���0�u�:�u�w�����8����I��QN����x��0�8�/�+��������p��T-�����<�u�`�{��8����Ӓ����X��ʶ�;�=�9�_�w�p����������G��U���0�!�4�u�?�$����W���l�C��\ʁ�u�:�%�;�6�8��������R��X�����0�"�0�u�%�>����ӓ��G��_�����7�3�0�_�w�p����Y����_��RN����� �0�u�:�?�1�W�������p��t������&�8�9�$�}����s�����*��ʘ�8�'�0�u�6�8����Ӕ��^F��RN�����3�!�0�7�1�8�W���Y����]��R��U���u�'�8�&�6�1�4�������F��E�����;�u��9��>����(ӕ��C
��d��X���0�"�;�u�8�5����Y����V��VN�����&�4�4�9�5�8�����Ʈ�T��^ �����u�4�6�9�#�2�}���TӒ��V��E��ʻ�#�'�=�9�w�2�W��� ӕ��C
�������7�3�0�{��}��������[��N�����x�"�;�u�8�0��������[��V�����9�u�0�1�1�2�W���Y������X�����0�0�4�u�6�-��ԜY����D��Q��U���;�u�#�'�%�)����������T�����u�&�3�;�$�4��ԜY��ƹK�`�����0�4�&� �1�/�����ƿ�R��t�����u�a�u�=�$�*�Ϫ�Ӌ��T�������u�x�u�"�w�(����Y����V��[�����<� �0�{��8����ӄ��U��@��U���0�d�u�4�'�8�W������F��V �����<�u�0�1�w�)��������]����ʶ�9� �4�<�9�<�ϩ��Ƥ�E� N�����&�u�x�u�1�8����������T�����<�u�<�<�?�.�Ͻ�����G��d��X���<�6�u�=�w�(����Y����W��NN�����1�u�=�u�2�2�ϼ�����D������u�-�'�u�6�-��ԜY����E��V��U���;�<�u�!�%�.�Ͻ�����G��N����u�4�%�0�w�;����ӑ��G��G�����x�"�0�u�#�;�����ƭ�P��B�����_�u�x�u�z�}�^ϊ�Y����V��C�����=�u�<�0�>�8���� Ӊ��G��T�� ���<�;�<�u�?�}����s�����T����� �<�&�u�?�}��������A��_��ʷ�u�:�3�2�%�9��������W����U���u��9��4�8�Y�ԜY����V��d�����>�_�u�0�>�W�W���Ӕ��Z��R
��]���%�0�9�|�#�8�}���Y���/��@�����;�'�&�!� �}�����Ơ�GF��C�����!�u�=�u�6�<��������R��V��U���u�x�u�&� �}����Ӆ��R��_�����u�r�{�u�w�}����,����V�������u�u�u�&�"�;�������	��R��H���e�|�_�u�w�}����Y���F��QN�����,�9�&�<�"�����H����[��N��U���u�&� �3�%�4���Y����P%��[������0�x�d�l�}�W���YӃ��Vl�N��U���u��9��4�8�:���
����P��U�����0�u�=�;�f�s�>�������R��C����� �4�<�;�]�}�W���Y����A��_��U���u�0�;�#�%�/�ϱ�Ӊ��@��RN��U���4��8�'�2�s�>���
ө��G	ǻN��U���x�;�!�6�:�8����Y����G��S��U���&�!�7�!�2�3��������TF��^�����u�u�u�u��;���������B �����}�y��3�2���������]ǻN��U���;�u�3�_�w�}�W���Y����F�R ����u�0�1�%�8�8��ԶY����A	��D�����0�9�|�u�5�:����Yӏ��A��Y	������8�9��<�}����Y���K�~��ʴ�0�<�u�0�2�}�ϩ��Ƹ�
��
��ʳ�:�u�:�!�2�9��������V��DN���ߊu�u�u�x�6�}�Ͻ�Ӓ��P
��EN�����<�=�e�&�]�}�W���ӕ��V��D�����_�u�u�u�w���������R��Y�����u�h�}�!�2�.�J���I����F�N���ߊu�u�u�u�z�.���� ����~��D!��U��� �1�;�#�%�?�W���
Ӓ��]F��@��U���0��&�!�>�}����W���F������;��9�,�>�(�2������@%��T-�����<� ��0�z�j�}���Y�Ʃ�WF��d��Uʰ�1�<�n�u�2�9��������9F�N�����u�0�0�y�#�8����Y����A��	��U���!�4�<�0�w�$� �������V��d��X���:�8�;�8�-�}��������W��Y	�����;�!�4�<�6�4�Ϫ�ӂ��RF��Q��ʴ�0�'�&�!�6�9�W��Y����Z��R
��ʸ�;�8�8�1�;�$�����Ʈ�U ��^ �����x��0�u��8�%���ӂ��@��C����� �3�'�<�w�1�Ϭ�
����\F�������:�u�:�8�;�2�������F��X���8�9��>�]�}����s���Z ��^�����2�}�4�%�2�1�^Ϫ����F�D;�����0��%�u�j�.��������9F�N��'���!�0��<�#�/�W��
����a��C>��ʭ�'�&�&�'�2�8�L���Y����a��C#��%���!�'��%�w�`��������c	��C��N���u�0�1�<�l�}����	����@��=N��U���=�:�
�u�%�>�3�������_��s��<���9�,�u�u�z�+����Ӎ��G��N=��ʾ�4�4�;�'��'�}���Y�˺�\	��VN�����u��&�!�2���������Vl�N����>�4�&� �1�/����
����V��MךU���x�=�:�
�w���������WF��V�� ���!�4�<�_�w�}�Z�������@"��V!��<ʦ�4�4� ��#�W�W���T����X9��D*������&�4�4�"���ԜY�ƈ�G��s�����;�<�,�"�%�s����=����G��[��]���|�u�u�u�0�3�������9F�N��U���8�4�4� �1�/�W�������R��B�����u�x�<�u�>�)����C����F�N�����4�'��/�w�}�J���=����]'��d��\���x�u�;�u�9�8��������F��\��H��u�u�u�%�%�}����s���F�D<�����u�u�u�u�w�}�W���Y����a��C#��%���!�'��%�{�}�W��Y���Q	��R��U���u�u��8�;�����Y���F�N��H���4�%�0�9�{�}�W���Y���F�C����&�1�9�2�4�}�W���Yӕ��C��Y�����<� ��2�#�`�W���	����V"��V�����<�=�y�u�z�4�Wϫ�
����WN��S�����_�u�u�u�w�����*����F�N��U���u�k�&� �1�/����Y���F�N��U���u�;�u�;�>�3�������\F��N��U���&�4�4�;�6�4�W���Y���F�
P��1�����9�1�w�}�W���Y���K�^ ��7���0�;�0�!�%�6����Y���F��s��<���u�u�u�u�w�}�W���D�ƿ�R��Y'�U���u�u�u�u�w�}�W������Z��S_�����
�}��_�w�}�W���=����]7�N��U���u�u�u�u�i�.�������F�N��U���u�u�x�u�9�}�����ލ�A��CF�����u�u�u�&�6�<�������F�N��U��u��!��1�(�!������F�N��Xʺ�!��:�0�9�8��������9F�N��U���!��!�u�w�}�W���Y���[�D*������!�y�u�w�}�W���Y���	��=�����m�'�g�
���}���Y���@"��V!��$���u�u�u�u�w�}�W���
����q��B��N���u�u�u�u�w�p�W���Y����V��v��1���>� �_�u�z�����Y����U��CN�����!�:�u�=�w�/����Ӣ��RF��E��[���&�4�4�4�>����Y����w��~ �����_�u��!��$�_���E�ƿ�R��Y'�Uʦ�4�4�'��g�}�Jϭ�����b]ǑN�����6�;�!�4�6�/����s�ƪ�AF��^ ��;���'�6�&�<�0�3���Y����G	�	�����0�u�u�x�w�<�Ͻ�����]F��X��U���>�4�4�;�%���������[��V�����0�{��u�6�}�����ƈ�G��C8���ߊu�u�x�3�%�<�Ϫ�ӕ��C
�������u�4�4�7�$�W�W���=����R
��v�����h�}�!�0�$�`�W�������|��V��]���|�n�_�u�w�p�6����Ƹ�VF��C�� ���!�u�'�8�#�8����Y����V��C�����4�4�4�'�.�s�W���>����\��^������,�o�u�w�;�ϴ��Ƨ�R��Y/��&���x�u�:�;�8�m��������F�N�����'��<�}�~�a�W�������|����Y���_�u�u�u��)�6���Q����F������3� ��<�f�7�L���YӃ����R��ʒ�;�'�6�;�#�<��������9F��Y
�����4�0��;�%�>��������A��dךU���0�4�0�'�4�1����s�ƪ�AF��X�����;�0�u�;�<�(�'���;����@K��S�����u�0�0�4�2�}�Wϭ�����R
��v����}�'�6�9�4�����Y���@5��E�����4�<�}�'�4�1�������9F������'�4�}�|��2�5�������KO�N��U��&�!�'��6�8�'���;����z��OG�U���&�0�1�1�%�.�6��� ���c��u�����0�|�i�u��<�6�������c�������1�0�&�;�>�8����P۶��P$��T�����n�u�u�&�4�(�6��� ����Z������h�u�:�=�%�}�I���^����F�D/�� ���'�,�}�|�k�}�������N��_��U��r�r�|�_�w�}�Z��������������<�2� �<�$�}�Wϙ�����V6��T;����u�u�3�'�>�4�W���Ӎ��^6��T�����;�!�u�0�2�<����Y�����X��U���6��6�'�4�3����Y�����X��U���'�!�;�=�>�}�J�ԜY���K��X��ʾ�:�3��8�9�)������ƹF�C�����
�u��"�$���������\��^��6ʦ�:�0�!�:�1���������@+����\���u�u�x�#�8�6�ϭ�����G%��Q�����:��<���.����
����U ��S�����<���<�f�W�W���Y�˺�\	��VN�����!�:�3�u��8��������C��d��U���x�#�:�>�6�.����)����e��SN������9�1�'�6�u�Z���)����_	��~ ���ߊu�u�u�x�?�2�(���*����c��RN������'�,�<�f�u��������]��d��U���x�#�:�>�6�.��������@/��D<�����'�&��'�.�4�F�������\��Y
��\���u�u�x�#�8�6�ϭ�����P6��D�����<�u��4�2�<��������N��X�����;�0�|�u�w�}�Z¨�������O�����&��!�&�?�.�6��� ۏ�c��u�����0�|�u�u�w�p��������a��v
����� �u��4��9��������ZO��E������1�-�_�w�}�W�������RF��V�����<�u��!��1����Q����9F�N��X���:�
�u��#��>ϭ�����J/��_��U���u�x�#�:�<�<��������@"��V/��$¼�d�_�u�u�w�p����&�ƿ�P��~ ����� ��'�,��p�^ǎ�����P��S�����u�u�x�=�8��W�������bF��T��4���,�}�x�|��2�5�������KOǻN��U���=�:�
�u��>����/������T������'�,�<��/��������V�N��U���#�:�>�4�$�>����������T������<�}�'�4�1�������F�N����>�4�&�6�"�����(ӕ��P��E��$¼�}�'�6�9�4�����s���F�A�����&�6� ��#�}�6�������A��~F��]���6�9�6��3�%�}���Y���E��\1����� ��!�u��>����8����bN��>�����6��1�-�]�}�W�������V��X�����u�;�<�,� �/�Y�������c��b ��U��_�u�u�w�}�����ơ�CF�N��U���u�>�4�4�9�/�$���Y���F��V������/�y�u�z�4�WϷ�������P��U���g�o�u�_�w�}�W���Y����@��t�����u�h�u�h�{�}�W���Y���K�^ �����0�;�u�u�w�}�Wϵ�����V��D�����k�<�d�u�w�}�W���Y����������_�u�u�u�w�2�ϳ�	��ƹF�N��U���0��&�!�w�}�W���Y���F�S����'�0�0�y�w�}�W���Y���F�N��U���u�u�x�u�9�W�W���Y���`��[�����u�u�u�u�w�}�W���Y����R��R-��Y���u�u�u�u�w�}�W���Y���F�N��Xʼ�u�u�u�u�w�}����
����A��Y��U���u�u�u�u�j�}�'�������V��CB��U���u�u�u�u�w�}�W���Y�����=N��U���u�u��"�$���������\��^��6���k�&�:�0�#�2��������A2��D#��]���|�u�u�u�w�p�W���s���F�N�����&��0�3�9�8�1�������pF������!�:�3��3�%���������B��U���u�x�<�u�w�}�W���Yӕ��_��T��8���&�;�u�u�w�}�W��Y����P%��[������0�u�u�w�}�W���Y���F�C���ߊu�u�u�u�w�����:����F�N��U���u�u�u�k�$�.�6�������Z��^G�U���u�u�u�u�w�}�W���T�ƥ�l�N��U���&�!�'��6�8����Y���F�N��H����4�0�4�>��������c��u�����0�|�u�u�z�4�W���Y���F��d�����&�u�u�u�w�}�W���Y���F��_��4���,�<�d�}�%�>����0����J�N��U���u�;�_�u�w�}�W���+����W��D��U���u�u�u�u�w�}�Iϭ�����W��D/�����x�|��:��2�������K�^ ��U���u�u�u�&�2�)��������G0��^
��U���u�h�u��6�8����8�����g��7���>�;�0�|�w�}�W����ƹF�N��U���-��6�=�$�����Y���F�S����&��'�,�>�u��������]��B��U���u�u�x�u�"�W�W���Y���@"��V'�����u�u�u�u�w�}�W���Y����w��a�����}�x�|�u�w�}�W���Y���F�N��Xʼ�u�u�u�u�w�}��������F�N��U���u�u�u�u�j�}�3���8����ZK��N��U���u�u�u�u�w�}�W���Y�����=N��U���u�u��!���W���Y���F�N��U���k�&�4�4�%����U���F�N��U���u�u�u�u�w�p�W���s���F�N�����1�'�&��#�}�W���Y���F������1�0�&�'�6�u�^ǎ�����P��S��Y���u�x�:�!�w�}�W���Yӕ��P��Y'��U���u�u�u�u�w�}�W��Y����F��E��]���|��:��8�6����P���F�C���ߊu�u�u�u�w��������F�N��U���u�u�u�k�$�>��������ZK��>�����6��1�-�{�}�W���T�ƥ�l�N��U���&�6� ��#�<����Y���F�N��H����6�8�4�>������Μ�\��X�����|�u�u�u�z�2����Y���F��v������9�u�u�w�}�W���Y���F��T��4���,�}�|��8���������F�N��U���u� �_�u�w�}�W���8����|��T��U���u�u�u�u�w�}�Iϭ�����A��fF��]���6�9�6��3�%�[���Y���K�X��U���u�u�u�&�4�(�8���Y���F�N��U���u�h�u��4�0��������ZO��E������1�-�y�w�}�W����ƹF�N��U���6�8� ��w�}�W���Y���F�S���� ��!�'�6���������\��Y
��\��u�u�x�u�"�W�W����ƫ�]��C�����4�0�'�6�9�)�L�ԜY���5��R�����3�;�9�4�4�0����Ӊ��C��d��U���u�:�<�0�#�<�W�������F��C�����'�a�u�<�$�2�ϱ�Y����R��Z�����u��<�u�$�.��������Vl�N�U���u�4�<� �w�8��������VF��G��ʥ�'�%�:�0�$�3�W����ƥ�W��N�����u�=�u�4�2�}�W��Y����V��V�����2�0�u�:�w�}��������	��^��Yʡ�<�u�0�1�w�2�ϳ�������^�����:�_�u�u�z�)�Ͻ�����Z��DN�� ���!�u�e�z�a�`�A������[��B��ʡ�0�4�&�9�#�}����Y����[ǻN��Xʷ�&�u�:�3�>�4�����ƭ�\��_�[���=�&�8�4�$�)�����Ơ�A��CN�����"�u�:�9�w�+�ϻ�	����F�C�� ���3�!�0�4�4�0����ӏ��H��@�U���{�b�{�u�1�*�W����Ƹ�Z��GN��U���u�0�!�%� �/����U���K�@�����z�e�`�8�/�}�$���ƭ�VF��Q�����<�2�4�4�w�5�W����ƪ�F��^�����=�u�6� �"�<��ԜY�����B�����<�=�4��b�m��������R��Y@ךU����6�8� ��1�ǎ�����P��S��U��&�6� ��;�9����Q����c��R�����<�&�}�'�4�1�������9F������ ���:��2�������F��T��:���'�4��>�"�����
����]��F�����:�>�;�0�~�6��������T��N�����u�|�_�u�w���������A	��[��<���-�u�h�&�4�(�8���������Z>�����<�2�;�!�~���������W�������!�0�2�=�f�9� ���Y����9F��Y
�����4�0��;�%�)�'���;����@]��Y
��!��