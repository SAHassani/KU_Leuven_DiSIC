-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:��:�>�8��!������r��X�?���u�8�0�8�9�p�W�������6��]��Oʅ��
�c�`�]�p�3���C����y��\�D���_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԑT�ί�T��N�����2�!��!�8�<�W�������]��t�����<�;�x�u�;�}����
Ӵ��V��Sd�U���<�;�9��$�/����
ӯ��V��[N�����4�<�;�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��ƴl�>�����o��<�u�>�8�����Ƹ�R��V��U���8�!�0�&�3�1����	������CN�����u�u�u�u�w��W�������Z	��y��U��� �'�1�!�w�5�W���T����_	��TN�����:�u�=�_�z�}�W���Y�Ɗ�R��Y�����6�9�6��'�W�Z��Y���F�=��ʦ�2�4�&�4�2�4����ӏ��G��N��6ʶ�&�{��0�>�-��������QǶN��U���u�u�&�1�6�9��������G��^�����:�;�6�0�w�2�Ͻ�����GF��:��ʦ�8�_�x�u�w�}�W�������@F��RN�����u�;�:�4�%�$�W������5�����߇x�x�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǑ[�����<�0�y�"�%�f�Wϫ�ӏ��VH��S1�����d�c�{�9�l�}��������]��E�����4�9�_�u�$�}����)����f��^�����{�9�n�u�"�8� ���W����A��~ �����9�n�u� �2�*����������d�����,��4�!�9�8��������X2��d"���ߊu�0�0�<��}�Wϵ�����@6��t����<�u�;�0�2�}����Y�Ƹ�T�
N����u��0�6�8�6��������]F��C��ʧ�;�0�g�!�w�}�J��B����\��=N��U���%�0�9�u�w�3��������l�N�����>�o�<�u�#�����B�����x�� ���&�o�<�u�#�����B���F��V�����0�;�o�<�w�)�(�����ƹF��s��'����1�0�&�1�.����Cӏ��@��[�����6�:�}�u�8�3���B���fT�=N��U���!��4��3�8����
����\��YN�����2�6�#�6�8�u�W������]�N��[�ߊu�u��4�2�3�W���ƿ�W9��P�����:�}�m�1� �)�W���Y����_�=N��U���4�0�;�u�m�4�W���&����P9��T��]��1�"�!�u�~�}�Zύ�@��ƓF�D*�����4�<�u�u�9�.��������F�D*�����e�o�<�u�#�����&����\� N�����u�|�u�x��e�F���Yӕ��G��~_��U���&�1�9�2�4�+����Q����\��XN�N���u�d�{�_�w�}�3���0����	F����*���<�
�0�!�%�l�W������]�N��M��u�u�&�4�6�3�F���ƿ�W9��P�����:�}�b�1� �)�W���Y����^�=d��Uʦ�6� ��!�6�4�W����ƿ�W9��P�����u��6�8�"��W����ƿ�W9��P�����:�}�`�1� �)�W���Y���`R�� d��Uʦ�6� ��!�f�g����
����\��h�����a�u�:�;�8�m�L���Tӵ��QǻN��4���8� ��u�w�(�W���&����P9��T��]���1�"�!�u�~�}�Z���M����F�D/�� ���!�d�o�:�#�.��������V��EF�U���;�:�e�|�w�p�W��W���WF��V�����%�'�6�9�4�	����B���P��R������u�3��6�)����	����q
��\:��&���<�_�u�x�w�/�����ƭ�A��C�����!�0�8�9�>��4Ϸ�	����2�������<�0�<�_�w�p��������WF����U���<� �u� �5�/����)�ƿ�C��C�����=�u���]�}����ӕ��G��E�����u�<�;�1�o�/����Q�ƨ�D��^����<�;�9�&�6�<����0���5��Y��M���4�
�}�u�8�3���B����Z��[N������'�,�;�m���������\��XN�N���&�2�4�u��)�%���8����@��Q��<���u�u�;�<�9�9�6��� �����Y��E��u�&�2�4�w���������T��N�����!�!�d�1� �)�W���s�ƿ�T������� ��<�;�3�}��������F��@ ��U���_�u�<�;�;�.����6����_��X��U���9�4�n�_�w�p����&����G��=N��X���:�
�<�0�3�W����s���6��\N��ʸ�9�<���������ƥ�G	��YN�����u�;�,�!�2�;����Y���X5��G��%���,�9�u�9�:�3�Ϸ�Y����R��NN�����0�6�;�0�#�9�W��Y����@��V��ʴ�:�1� �;�4�.����?���F��V�������i�u�$�:����=����]/�������&�4�4�;�g�t�}���=����A��~ ��I���&�2�0�}��)�>���Pߕ��]��D*�����e�|�_�u��<��������[�B �����}��4�0�9�t��������@6��D��E���_�u��!��<�6�������U��~ ��U��}�;�<�;�3�.��������W��D!�����|� �&�2�2�u�3���+����W��D�����e�|�_�u�z�}��������[��G�����!�u�'�6�$�4��������l�C�����2�;�'�!�w�1��������\F��A�����7�9�!�u�9�)�Ͻ��ƻ�����U���=�u�x�u�6�8�}���T����X9��q�����0�%�'�6�;�>�#���Y����[	��h��0���!� ��&�#������ο�])��G��3���u�x�#�:�<�<��������_��X1�����;�&�4�6�9�?����s���E��\1�����&�u��4�2�/����Q����C
��g�����u�u�u�:�9�2�G�ԜY�˺�\	��VN�����0�1�1�'�$�����0�ƿ�R��R�����&��3�0��u�$�������A%��[��U���:�;�:�e�]�}�Z�������@"��V'�����u�:�7�:�2�3��������_��=N��X���:�
�u��#��>ϭ�����A��Y'��&���9�&�0��4�8�Z������\F��=N��X���:�
�u��#��&ϭ�����A��Y?��&���9�&�0��4�8�Z������\F��=N��X���:�
�u��4�0��������r��Z!��#���1�:�9�u�z�+����ӕ��P��B����� ��!��0�8�_�������c��N��U���u�:�;�:�g�W�W�������RF��T��:���u��6�8�"�����ۍ��^��D>��6���0�x�d�1� �)�W���YӠ��P��C��%����:�>�:�/�}���� ӑ��XH��V�����%�'�6�9�4�	����-��ƹF��R �����4�u�_�u�w�}�$�������A%��[��Kʾ�4�%�0��%�$���Y����]F��Y�����4�2�u�u�8�o�M���s���F��A������6�:�u�i�6��������R��EG��X���;�u�;�0�2�}����Y�Ƹ�U�
N�U���%�'�u�4�w�W�W���Y����_��\N��U���u�u�u�u�w�c�$�������l�N��:����>�u�u�w�}�W���Y���X��A�����u�u�u�&�9�(����?���F�N��U��u�:�7�:�2�3��������u ��d��U���&�4�6�;�5�8�W���Y���F�
P�����:�0�;�&�6�>�������9F�N��%���0�u�u�u�w�}�W���Y���F��_��4���,�;�>�4�'�8�'��� ����F��S�����|�_�u�u�w�����/����F�N��U���u�k�!�
�8�1����=����]0��^
�����u�u��!��<�6�������U��~ ��Kʦ�4�4�0�1�3�/��������]N��V�����'�,�9�u�w�}�������9F�N��1�����u�u�w�}�W���Y���F��V�������>�4�'�8�'��� ����F��S�����|�_�u�u�w�����(���F�N��U���u�k�&�4�6�/����(ۍ��^��D>��6���0�x�d�1� �)�W���s���F��T��:���4�<�u�u�w�}�W���Gӕ��P��B�����:�9�_�u�w�}�6�������F�N��U���u�u�k�&�4�(�8���*����WN��V�����'�,�9�u�w�}�������9F�N��4���8� ��u�w�}�W���Y���F��T��:����2�0�}��0��������_�_�����:�e�|�_�w�p�6����ƃ�G��Dd����� ��!�4�>�}�K�������_	��TF������!�4�<��2�^�ԜY����F��C'�U��&�1�9�2�4�+����Q����F��C'�����}�|�n�u�$�>�������[��C
�����
�0�!�'�$�>��������]��G�����6�8� ��}�K�������T��A������6�8� ��4����H����[��\=������'�,�9�w�}�W����Σ�[��S�R��n�u�&�6�"����Y����G��X	��*���!�'�&�6�"���������O�@��U���8�9�&�0��>���KӃ��VF��C����u�e�|�_�2�9�%���s