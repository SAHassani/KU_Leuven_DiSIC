-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��G@�����u� �=�'�w�<�W�������\��t�����4�1��0�?�3�3���s����A��Y��%���0�!�u��2�h�Cڌ�T�ƈ�G��N�����e�e�x�_�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�TG��E���%�'�2�#������ƅ�@��Z��ʖ�'�:�4�<�9�p�W���Y����G��R�����x�u�4�<�9�1�>�������G��Y������3�'�4�>�3�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=C�X��� �%�&�o�z�}�W���Ӣ����[חX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�W�����ƥ�V��X�����&�u�0�0�$�9��������H��[UךU���u�0�0�;�:�/����݇��l�B�����{�>�� �>�4����
�ȭ�_]Ǒg������2�&�u�$�W�W��-����P��C����� �%�'�u�"�)����
����V��R�����{�u�!�%�w�4����A����J9��^�����u�u�4� �6�}����E���\ ��^	����u�:�;�:�g�f�Z���H����9F��B �����!�
�9�`��}�W���������B�����9�2�6�#�4�2�L�������Z	��C����}�u�u�;�2�8�^Ϭ�����@��[�����6�:�n�u�1�3����Y����^�����<�!�2�'�w�8��������V��N�����:�u�4�<�"�}����Y�ƥ�G��EG�����;�<�!�2�%�W�W���������[��U­�o�<�!�2�%�f�������]���� ���<�!�2�'�]�}��������^��R���� �&�2�0�l�$�MϷ�����O��R��ʼ�!�2�'�_�w�(����ӕ��_
��F��U���u�;�<�;�3�}����ӏ��V��d�����!�:�u�:�e�8��������Z��P��U��� �;�<�!�0�/�}��Ӷ��w��=d�����0�7�1�u�<��Ϸ�s����F��^�����9�`�}�u�w�3����PӔ��F��D�����6�#�6�:�w�.�Wϼ���ƹF��R��ʦ�1�9�2�6�!�>��������Z��SF��U���|�_�u�;�w�(����Ӓ��`
��dךU���6�<�;�!��1�O���Y�ƥ�G��EG�����;�&�1�9�0�>�����ƥ�9F��R	�����u�0� �;�$�9��������G	��C�����;�1��u�o�t�}����ƪ�]��X �����d�n�_�u�"�>��������F�OB��U���;�0�0�|�%�)��������AF��=N�����_�u�u�3�/�a�Ϫ����F�E�����n�u�u�0�$�W�W���Y����A��d��Uʰ�1�<�n�u�2�9��������^��Z�����3�;�!�:�w�<����Y۞�JF��^ �����u�0� �;�>�)�������Q��Yd��Uʼ�u�u�u�u�?�3�W���YӔ��F��OUךU���9�0�u�u�w�/����Y��ƹF��Y
���ߊu�;�u� �4�4�ϳ�����lǻ�����;�&�4�9�%�u�MϷ�����F��N�����0�|�'�!�%�}�����ƥ�9F��R	�����u�&�0�!�.�5����Y��ƹF��R�����;�<�;�1�%�3�Ϸ�Y����_��RN��U���6�8�4�0�w�2��������ADǻN�����<�,�0�'�%�W�W���������[��]���:�<�!�2�%�$�^�ԜY����U��C��U���9�0�n�_�w�(����ӕ��_
��F��U���<�;�1�u�w�}��������V��YN�����'�<�_�u�2�4�}���Y����A������f�_�u�u�2�2��������V��V ��U���!�:�9�'�2�)�W�������A��C��ʼ�!�2�'�_�w�}��������A��d��Uʧ�!�'�u�8�;�8�_�������V��B��N���0�1�3�;�#�2�W�������9l�Q�����u�8�9�0�w�%�W���Y����T��N�����u�;�0�0�w�.�Wϼ���ƹF��D��ʭ�=�2�u�u�e�<�ϧ�����F��=N��U���:�!�w�;�>�3�Ϭ�����@F��XN�����!�u�0� �9�4�P�������R��YN�����'�_�u�u�2�8��������l�N�����u�8�9�0��2��������J��h�����}�|�n�u�2�9��������@��[�����x�u�:�g�2�.�W�������_	��v��X���:�u�'�k�w�3�W�������F��EN����_�u�x��0�u��������A�^ �����>�� �<�>�4����Y����A��A�����'�8�e�!�w�3���� ���K��_����� �&�'�6�w�}�Ϫ�Ӕ��F
��X����%�&�!�#�w�/�^����ƭ�'��T��D���x�u�=�;��:�_���T���K��:�����1�!�<�u�2�<��������GF��^�� ���<�;�=�;�;�.�W��Y����r��S��U���0�"�!�u�9�8�������F��Y�����:�g�0�&��/�W�������AO��R��ʼ�!�2�'�<�]�}�W�������4��B�����u�;�0�0�l�}���������v��H��!�0�_�u�w�}��������	[�d��Uʰ�&�_�u�u�w�8��������*��F�����u�n�u�u�2�9���Y����V��YN������9�_�u�9�}��������9��>��1���_