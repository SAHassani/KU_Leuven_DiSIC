-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:��:�>�8�s��ԑTӧ��[	��$��ʔ�8�'�4�u�9�}����:����]	ǶN�����4�u�'�?�4�g�'���&����al�*�����l��9�u�g�l�Z�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���6�u�e�d��-����Ө��Z	��[N�����8�;�&��%�2�������r
��e�����0�0�#�1�z�}��������]��B�����;�0�;�9��;������ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�x�u�"�-���Y���� ��RN�����&�4�%�:�2�.��������U	��C�����!�:�4�_�z�}�W���Y����]��G�����u�!�!�>�$�4�W���Ӊ��G��d�����>�1�8�<�y�}���Y���F�N�����:�0�u�=�w�<�Ϫ�Y����|��t�����<�u�=�6�w�.��������WF��R���߇x�u�u�u�w�}��������p
��N��ʱ�2�!�9�&�0�<�W�������]��DN�����;�!�0��2����Y���F�N�����u�;�u�=�9�)�ϱ�����W�������&�0�'�1�5�>�W�������R��R-�����u�u�u�u�w�9����W���K�N��U���u��0�6�8�6����ӏ��Z��R�����4�,��0��6�����Ƹ�V��V��X���u�u�u�u�w�2�W���ӵ��C
��[�X�߇x�u�u�u�w�}��������C
��g�����u�;�<�4�2�5� ϳ��ƿ�^��DN�����;�<�,�x�w�}�W���Y�ƾ�P��R��ʡ�0�&�4�4�9�r�W������@"��V'��Z���'�u�4�&�3�p�W���Y���F��@ �����u�;�4�&�9�1�W���Y����F��T�����;�u�;�!�2�<�������F�N��U���4�&�1�:�w�}��������|��T��ʶ�6�0�u�:�w�5�Ϭ�����K�N��U���u��%�!�6�-��������VF��R
�����0�&�4�9�%�)����Ӄ��R
��Xd�U���u�u�u�u��8�4�������\�CחX���u�u�u�u��4�W�������G��DN�����6�9� �4�>�3���� Ӓ��VF��V�����0�x�u�u�w�}�W���
����@H�u��ʺ�u��4�0�w�)� ���Y������T�����=�u�<�!�%�2����s���F�N��U���6�8� ���2����Y������A��ʢ�0�u��6�:�(�!���Ӈ��V��N���߇x�u�u�u�w�}����Y����[��R
�����!�0�&�<�#�/��������JF��D�����&�4�4�;�6�4�}��Y���F���ʣ�9�1�1�!�w�4�W�������XF��T��U���0�u�;�&�6�<����WӲ����VחX���u�u�u�u�$�2����ӏ��_��Y��U���!�0��7��
�1���Y����A��=C�X���u�u�u�u�w�5�W����ƨ�G��R�����0�&�u�;�w�5��������[��
�����;�u�<�0�>�8�Z���Y���F�S��ʦ�'�6� �0�y�	�ϲ�����V��E�����;�<�0�"�.�)�W����ƭ�_F��Rd�U���u�u�u�u�6�5�[Ͽ�Ӂ����ZN��U���6�u�=�u��}����Y����[��V�����u�&�!�_�z�}�W���Y����V
���������<�u�?�}�!Ϛ�����F��V�����u�=� �1�%�<�Ϫ��ơ�W��=C�U���u�u�u�c��8�4�������@F��C�����6�;�7�0�w�3����ӑ��W��s��<����8�&�_�z�}�W���Y����VF��[����>�#�'�9�4�����Y����V��X�����u�=�u�0�#�2�W���Y����GǶN��U���u�u�<�u�?�}��������W	��^ �X���u�u�u�u�w�2�ϭ�����e��SN��ʦ�4�4�0�1�3�/��������]F��RN�����0�%�6�0�w�2�Z���Y���F�U�����4�<�;�1� �)�W�������_�u��U���!�<�u�<�9�1�W���Y����	��=C�U���u�u�u�6�4�8�����ƿ�R��Y'��U���u�!�<�u�8�}��������\F��A��U���'�9�_�x�w�}�W���YӅ��_��X�����u�;�!�0��}������ƴl�N��U���u�u�:�u��0��������_�\����4�0�1�1�%�.�8�������P	��V��U���<�!�2�'�z�}�W���Y���\ ��R�����!�u�2�:�2�)�ϸ�����R��R��ʡ�0�&�<�!�%�:����
�Ƙ�Z��Dd�U���u�u�u�u�2�9�ϼ�������*��ʶ�8�&�<�u�%�(�ϱ�Y����C
��g�����y�"�<�=�:�<���Y���F�N�����1�!�u�4�w�8�����Ƹ��������&�u�#�;� �8�W����Ƣ�GF��CN�����u�:�_�x�w�}�W���YӒ����E��U���6�9�!�:�y�����
����a��v
�����3�&�!�;�!�1�������D�^����u�u�u�u�w�<����I��ƴF�N��U���u�e�u�k��8��������GF��C�]���8�;�u�u�1�)�ϲ�
�ƺ�_��S��Y���u�u�u�u�w�}�W���Y�ƥ�P
��^ �����1�!�u�=�9�.��������WF��D�����x�u�u�u�w�}�W���H���f��C�����;�u�0�0�#�9���Q����V��N��U���u�4�!�#�;�9����U���F�N��U���u�u�u�<�4�(��������R��@��U���!���9�3�<����
��ƴF�N��U���u�d�u�k��8����������R�����{�x�u�u�w�}�W���Y���F��^��ʻ�!�4�#�9�3�2����W���K�N��U���u�=�&�8�3�1�W���������R�����!�u�0�!�"�}����Y�ƀ�u��
�����u�0�0�_�z�}�W���Y����V��R��[���_�x�u�u�w�}�Wϊ�Ӗ��V
��RN�����!�'� �=�#�4�W�������@l�N��U���u�u�:�;��u�E���M���O��x�����>�4�!�'�w�}�W���	����XF��T��[���_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�Զ����A��R��U���>�_�u�&�w�8��������Z��X����_�u�&�u�2�8��������G��[�Uʠ�0�"�'�{�<��"�������w��V�����&�u�:�>��:������ƹ����ą�2�'�6��#�/�Y���B���G��(�����!�'��:��2����Y��ƹ��R��]���u�>�4�%�2���������Z��Y�����4�2�u�u�8�o�M���B�����R�����4�!�'�o�>�}�����ƾ�]��N��U���h�f�n�u�'�/�_���Yӵ��C
��[��U���&�1�9�2�4�W�W�������XF��^ �����:�<�n�u�w�.����	����@F��^ �����4�n�_�u�w���������	F�������n�u�u�&�?�.�W���Ɯ�R��CF�����0��'�,�;�p�W������]�N��L��_�u�u��#��!�������]F��X���ߊu�u��!��<�6�������U��~ ��U��� �&�2�0�e�/����Q����C
��g�����x�u�:�;�8�m�L��Y���9F�������o�<�u�>�3��������GN��V�����'�,�9�x�w�2����I���F��@�U���&�4�4�;�w�}�ύ�����'��V��]���8�9�&�0��>�������\F��N�U��{�_�u�u�$�>��������WF��X�����0�;�_�u�w��������	��*�����
�}��8�;�.���������Y��E��x�u�a�{�]�}�W�������G7���U���4� �
�}��0��������_�
�����e�|�u�x��k�@��Ӡ��P��C��%����:�>�:�l�W��������A��c"��ʓ�4�!�;�0�'�/����������N�U���u� �7�'�8�}����
����3��C�����1�7�u�4�6�1�W�������^��^ ��U���u��9�%�6�8��������G��B�����4�<�;�x�4�(��������C��T���ߊu�x�>� ��2��������G�-�����}��9�%�6�8��������G��x�����>�4�!�'�]�}��������}��E�����2�;�!�u�w�<����s���F�N��U���u�u�u�u�w�}�W���D�Χ�\
��_��3���0��;�!�w�}�8�������u��X��U���z�>�#�'�;�>�1�����ƹK�c�����!�u�3�!�2�;��������D	��R�����4�u�4�0�"�1�W�������l�C��<���!�,�6�=�$�6��������R��EN��Dʓ�&�4�1�:�"�-����ӎ��9F�N�����9�6��6�8�}�1��4����W��^�����1�&�'�7�3�4�W���Y����V��N�U���!� �0�u�?�.�������F��P ��U���!���;�w�}��������G	��\!�����6��6�:�w�2����I����N��_��U��3�9�0�n�w�.����Y����F��Y��U���9�4��6�8�u�8�������u��X�����:�e�u�h��)����D�ƪ�_��d�����4�u��!�"�����Y����V��R��¾�#�'�9�6��>���Y����G	�N�Uº�=�'�u�k�1�1���s�ƿ�T�������4�9��%�w�}�������� ��D�Uʦ�2�4�u��#��!�������\��X�����h�3�9�0�]�}����ӕ��R��^��Oʅ�4�0�!�>�6�-��������VK��S�����|�o�u�:�?�/�J�������@F�I�\��x�u�g�{�]�}����ӕ��G��V
�����&�3�&�!�9�4���,����]��v�����>�4�%�0��/����T�ƨ�D��^��O���:�=�'�h�w�2����Y���A�N�U��g�u�&�2�6�}�3���0����V/�=�����m�'�4�
������
����J��_�����:�e�u�h��)����D����G��DN��R��|�u�x��o�l�Wϭ�����@"��V'�����u�u�<�;�3�e����&�Χ�R��R�����9�x�u�:�9�2�G���D�Σ�[��S�]���0�&�h�r�p�t�W��*���9lǻ�����:�4�6�;�5�8�Mϼ�����\�Q���ߊu�<�;�9�8�<��������	F��X����u�4�&�n�]�}����Ӊ��G��V
�����&�3�&�!�9�g�"�������r��N1�����%�0��'�.�1�Z�������V�S�����'�h�u�:�?�/�W���^���F�;�G���&�2�4�u��<���)����l��d�����0��6�0�f�9� ���Y���F��C����}�!�0�&�j�}�G���B���fU��d�����4�u��!���Mύ�����'��V��]���8�9�&�0��>�������\F��T��]���0�&�h�u�8�5����G���]�N��M��u�&�2�4�w�����(����Z��S_�����
�}��8�;�.���������Y��E���h�}�!�0�$�`�WǱ�����X�G�U����m�d�u�$�:����=����]5��^��U���<�;�1�d�w�2����I����N��_��U��e�|�u�x��e�F���
����_F��V�����<�9�u�u�>�3���Y����G	�N�Uº�=�'�u�k�g�t�W��*���9l�D������4�!�4�4�<��������]F������u�&�2�4�w�����/����t��N�����;�o�u�4�$�f�}�������	��T�� ���9�1�u�:�;�<�W������lǻ�����:�6� ��#�<����	����Q	��R��O���4�&�n�u�$�:����8����|��^��U���4�4� �
������
����J��_�����:�e�u�h��)����D����G��DN��R��|�_�u�<�9�1��������c��fN�1����!�!�>�6�-��������VK��S�����|�o�u�:�?�/�W���Q����A�	I�\��_�u�<�;�;�.����6����_��T��U���
�:�<�u�j�z�P�ԜY����R
��v������9�u�u�6�<����Q����C
��g�����x�u�:�;�8�m�W��Q����A�	N�����&�h�r�r�~�}�Zύ�O��ƹ��Y����� ��!�6��g�3���6������Z������6�0�d�3�*����P���	��R��H���:�=�'�u�i�m�^��T�Ɵ�H��=N�����9�:�4�4�9�3�������]��[�����d�>�#�'�;�>�1����Ϩ�D��^��O���:�=�'�u�i�z�P��Yӕ��]��X=�����;�o� �&�0�8�_���K����N��A������6�:�|�8�3���B��ƹ��E�����4�
�4�:�#�}�������R��^��ʸ�-�3�;� �w�;��������PF��D�����&�w�w�_�w�p�W���
�ƿ�T��DN�����u�>�0�w�6�)����Ӓ��V��E�����!�0�u�:�p�}��ԜY����F��SN������f�&�u��8�ϰ�����\F����ʹ�2�6�%�!�w�8� ���Y����F�=�����9�u�;�u�!�/��������@F��EN�����{�u�4�!�>�(�ϵ�����@��Y	�Uʴ�!�<� �0�<�8�W�������v��[��U���;�9�<�u�#�(�U�ԜY����Z��RN�����3�:�4�4�2�9����
����@��YN����4�u�&�w�%�8�L�������Q����ʺ�u��!���1���
����_F��L�� ���_�u�!�'�5�)�W���	Ӊ��\6��D��U���;�9�<�u�#�(�U�ԜY����Z��RN�����3�:�4�4�9�}�W�������@F��E��N���4�!�<� �2�6����Ӊ��G��fN����4�u�&�w�%�8�L�������Q����ʺ�u��6�8�"�����Cӕ��]��^�����w�_�u�!�%�?��������UF��T��:���u�u�<�;�;�4�Wͪ�����F��C�� ���>�0�u�3�$�>��������@��V�����'�0�n�_�w�p�#���ӕ��]����ʴ�w�0�%�u�#�/����Y����]��RN�����=�,�1�;�#�:����T�ƿ�P����ʆ��g�{�u�?�/�W����Ƹ���VN��U���<�u�4�=�5�)������ƹK�x��6���4�1��8�;��Ϻ����� �������_�u�!�'�5�)�W���	Ӊ��@'��B�����<��9�u�>�3�Ϸ�Yђ��VD��N����� �0�>�0�w�;����������N�����u�&�w�'�2�f�WϿ�����G��R������6�8� ��1�Mϭ�����Z�C��W�ߠu�x�u�;�"�8����Y����@�������0�&�2�4�w�2��������^��Z�����<�=���w�2�W�����ƹ��E�����0�%�:�u��-�����ƿ�T����W���0�n�u�4�#�4��������\ ��s��<���;�o�&�2�6�}�������9F��C�����u�0�%�:�w�����*������Y�����!� �w�_�w�p��������@��Cd�����4�u��6�:�(�>�������G9��\=������'�,�9�z�}�������9F��^	��ʺ�6� ��!�m���������`��[�����6�0�d�1� �)�W���s�ƿ�T������� �!�4�<�m�?�������K��X�����;�_�7�2�9�}�Z�������G��^ ��ʦ�2�4�&�<�w�5�W���	����XF��Z��U���:�0�!�0�w�/�W���Ӓ��F���U���'�9�u�:�6�3�Wϊ��ƥ���RN��U��� �0�!�0�2�4�W���ފ��ZǻC����u�0�"�0�w�5�W�������U	��C�����u�%�:�0�$�����:���F��P��U���<�u�<�<�0�8��������p
�������u�u�&�4�4�3�������F�N�U���9��4�9�l�}�W���
����z��[�����u�u�u�i�w�����/����l�N�����4�0�1�1�%�.�8�������Z��N��U���h�&�4�4�2�9����
����@��YUךU���u��4�0�>�8�W���Y���F�
N�����n�u�u�u�$�<��������F�N��U��u��!���W�W���Y����R/��^��U���u�u�u�u�j�.������ƹF��Y
���ߊu�;�u�'�4�.�L�ԜY����R����U��� �u�<�;�;�}�Ϫ�ө��A%��
�����u��<�u�$�9����Ӄ��F��N�U���'�u�&�4�9�p����Y������@��U���u�:�4�;�1�/������ƹK�c��U���:�1�&�!�8�}����?������XN�����&�4�1� �;�}��������V��_��U���u�'�!�6�$�)�Ϭ�
�ƣ��������;�!�<�u������Y����R��T�����u�&�0�!�8�W�W���Ƹ�VF��(��4ʱ�4�'�8�'�$�)�}�������@N��R���ߊu�0�<�_�w�}�Ϭ�
����V��!�����|�!�0�_�w�}�W�������Q
��S��6����4�9��'�f�W���YӉ��G��a����u��!���1�������F�X>�����h�&�=�&��-�L���Y����w��e��4���0�&�3�&�#�3�K���=����V��S
�����3�0���'�f�W���YӉ��G��~N�U���!���%��W�W���Y����R/��R�����4�;�<�0�l�}�Wϻ�ӏ��9F��Y
�����&�n�_�u�z�����Y����\/��B�����<�;�9�!�6�}����Y����|��t��3���"�0�u�:�$�0��ԜY����R��Q��U���u�4�%�0�;�}��������A��RN��ʺ� �%�!�,�4�.����Y������[ךU���!�0��0��6�����Ɗ�@F��R ��ʹ�!�=�!�0�3�)�W�������G��X�� ���4�%�0�9�]�}�ZϺ�����u ��P�����:�'�6�9�y�}�Z¨�����)��E�����2�,�6�:�9�8�}���T����X9��\!�����6��6�:�w���������P��=N��X���:�
�u��"�)��������U��=N��X���:�
�u��$�)���������X��U���0�9�u�4�'�8��ԜY�˺�\	��VN�����u���!�"�����Tސ��\��!�����u�#�'�9�]�}�Z�������\%��Y��&���� �!�u�z�+����Ӊ��F��V��U���;�� �!�6�4�}���T����X9��X,������2��-�w�-����6����_	��^ �����:�;�0�-�w�3��������|��T������;�� �#�/�_���P�����R��U���u�_�u�u�w���������P��S����'�9�6��4�2�[���Tӏ����R	��U��f�u�u�u�<�2��������F�
P��F���u�u�u�u�w�}�W��Y���@��Y	��H���e�_�u�u�8�)����Q���F��e�����u�u�u�u�j�}����U���F�N��X���;�u�:�9�6�W�W���Y����p
��N��U���u�k��8�;�����Y���K�^ �����9�2�6�u�w�}�������F�N��H�����!� ��.�W���Y����]F��X�����h�!� �_�w�}�W�������F�N��U���0��>�w�}�W���Y���Z�D�����6�u�u�u�8�2����Y���F�
P��&���� �!�u�w�}�W������]��Y�����9�&�d�>�!�/����?����AO��=N��U���� �!�4�>�}�W���D�ƣ�J��X��#���1�u�x�u�"�}�������F�X,������2��-�w�c����P���F�N��U���:�!�7�:�2�3�}���TӶ��V
��RN��ʦ�;�u�<�;�;�}�ϳ��Ƹ�^�������!�u�0�!�w����� ����@F��G�����u�x�u��2�>��������M������u��!� ��3�W�������P��T��U���9�&�_�u�z���������p	��CN��U���u�,�6�1�#�}��������p
��R
��U���0�<�!�9�w�;�����ƪ�A��N�U���0�<�u� �$�<��������\�������'�u�0� �2�2��������R
�������u�;�u�;�.�>����T�ƣ�\�������&�;�{�u�'�2����6����_�N�����u�u�<�u�>�4�����΃�V��\G�����u�u�u�x�w�<�����ƥ�C��D�����4�0�'�2�$�8��������Z��_�����0�9�u�:�6�3�W���Y���R��C��U���!�0��0��6��������[��Z��ʚ�0��>�&�0�<�ϩ��ƫ�Gl�N��X���=�<�u�0�w�<�����Ƹ�VF��T��U���0�:�u�#�%�1�W����ƭ�A��Y	ךU���u�x�0�2�w�;�$�����������ʡ�0�'�#�9�2�6��������R��EN�����{�u�u�u�z�}��������_��g-����� �0�u�;�8�<�����ƿ�T��������;�� �#�<�W���s���F������;�u��!������
����@F��X��U���9�&�!�u�%�)�W�������c��N�����u�u�x�<�#�}��������V��N@ךU���u�x��u�!�4�W�������]��V�����4�u�:�0�#�<�W���ӑ��^��������9�1�"�#�W�W���Y����z��C=�����u�u�x�u�8�8����Y����`��[��ʱ�8�<�u�0�$�8��������\��B�����!�0�4�6�:�1����Y���K�@�����!�0�:�!�"�}�����ƹ�Z��x�� ���;�{�u�u�w�p�}���Y���.��RN��U���<�2�4�u�8�4��������[	��C��&���u�<�;�9�w�/�W�������l�N��X���u�u�u�u�w�}�W���&����l9��N��U���u�
�
�
��}�W���Y�Ɠ�l9��h1ךU���u�x�u�4�'�8����Yӹ��F�N��	���
�
�
�u�w�}�WϢ�&����l9��N��U���
�
�
�
�]�}�W���T���F�N��U���u�
�u�u��}�Wρ�Y����lF�1��U���
�u�u�
�w�}�(���Y��ƹF�C�U���'�9�u�u�w�����&���O9��N��*���)�
�u�)��}����YӚ��OF��h1��U���_�u�u�u�z�}�W���Y���F�N��*���
�
�
�
���(���&����l9��h1��*���
�
�
�
���(�ԜY���K�X-�����9�1�u�
�]�}�W���T���F�N��&���� �!�u�w�!�W��������N��U��u�u�d�u�w�o�W���I�ư�W�KN��Uʩ�u�u�u�x�w�}�W���Y���F�N��U���
�
�u�u�w�}�W���Y����lF�N��U���u�
�
�
�w�}�W��YӉ��C��N ��E���
�
�
�)�w�}����&����l9��N��U���
�
�
�
��}�W���&����9F�N��X���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�
���W���Y���F��h1�����u�u�x�u��-����ێ��[O��h1��*���
�
�
�
���(���Y�ư�l9��h1��*���u�u�)�
��W�W���Y���F�N��U���u�u�
�
���(���&����9F�N��X����9��4�;�}�(���Y���F�N��U���
�
�
�
���(���&����l9��h1��*���
�_�u�u�w�p�W���Y���F�N��U���u�u�u�u�w�}�W���Y����l9��h1��*���
�
�_�u�w�}�Z���:����]��RN��*���
�
�
�
���(���&����OF�N��U���u�u�u�)���(���&���F�C��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�
�
�]�}�W���T�ƣ�G��t��2���u�
�
�
���(���&����l9��KN��Uʩ�
�
�
�
���(���&����ll�N��X���u�u�u�u�w�}�W���Y���9��h1��U���u�u�u�u���W���Y���F�h1��*���u�u�x�u�8�<���� ���F��d>��	���u�)�
�
���(���Y����l9��h1��*���u�u�u�
���W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��*���
�u�u�u�w�}�Wρ�&��ƹF�C�U���!���;��4����Y����l9��h1��*���
�
�u�u�w��(���&����OF�N��*���_�u�u�u�z�}�W���T���F�N��U���u�u�u�u�w��(���&����F�N��*���
�
�
�u�w�}�(���&����l9ǻN��U���u��!���3�_���Kӵ��l�N��U���u�
�
�
�w�}�W���Y�ư�l9��Kd��U���x�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�(���&����lF�N��*���
�
�
�
�w�}�W��YӉ��G��d��]���=�u�u����(���&����l9��N��U���u�u�
�
��W�W���Y��ƹF�C�U���u�u�u�u�w�}�W���&����l9��h1��*���u�u�x�u�$�<��������l9��N��U���u�u�u�u�+��(���&����l9��h1��*���
�
�
�
���W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��*���
�
�
�
���(���Y���F��s��<���9�1�
�
���(���&����l9��h1��*���u�u�u�u�w�}�W���&����l9��h1ךU���u�x�u�u�w�p�Wϱ�����e��S)�����u�u�x�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���&����F�N�U���u�u�u�u�f��4���&����l9��h1��*���
�
�)�u�w�!�(���&����l9��h1��*���
�u�u�u�z�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y�Ɠ�l9��h1��*���u�u�x�u�w�}�W���Y����c%��h1��*���
�
�
�
���(���Y���F���*���
�
�
�
���W���Y���F�N�U�������}�w�]���S���L�D��_�������}�w�]���S���L�D��_����u�u�u�z�}�W���Y���F�N��*���u�u�u�u�w�}�W���&���F�N��Uʊ�
�
�u�u�w�p�Wϱ�����`��^��	���u�)�
�
���(���Y����l9��h1��*���u�u�u�
���(���&���F�N��U���u�u�u�u�w�}�W���Y���F��h1��U���u�u�u�u���(���Y���F�1��*�ߊu�u�u�x�w�����*����[��1��*���
�
�u�u�w��(���&����OF�N��*���
�
�
�)�w�}�W��Y���F�N��U���u�u�u�u�w�}�W���&���F�C����� ��!�4�>�}�W���&����l9��N��	���
�
�
�
���(���&����l9��h1��*���u�u�u�x�w�}�W���Y���F�N��U���u�u�u�u�w�}�(���&����l9��h1��U���u�x�u�:�4�(�8�������Z��h1��*���
�
�
�)�w�}�W���Y���F��h1��*���
�
�
�
��}�W���T���F�N��U���u�u�
�
���W���Y���l9��h1��U���u�u�u�
���(�ԜY���K�d�����>�u�u�
�w�}�W�������l9��KN��U���u�
�
�
��!�W���Y�ư�l9��h1�����u�u��!������DӉ��G��d��]���!���;�p�4�������\F��=N��U���u�u�u�u�w�}�QǱ� ����F��V��U���u�:�,�6�8�3�W���*����V��E-�����n�u�u�u�8�3�������	��G�����:�;� ��9�z����Hӂ��]��GךU���u�u�u�u�w�}�W�������p	��C8�����;�u��;��(���Q���9F�N��1�����1�-�k�}�$���:����l�N�����%�!�,�6�k�}�8�������PN��B�����6�=�2�x�w�2����I���F�N��U���u�u�u�s�8�$��������Z��Y
��&���� �!�h�<�+��������G	��N�N���u�0�1�<�l�}����	����@��N������9��!�w�}�W��Y����P#��U�����:�;� ��9�u�>���������_G�Uʺ�4�4�;�4�>�����Y���\"��V'�����u�;�u��#��$���Q����F��Y�����n�u�x�u�8�.�����Ƹ�VF��[�����9�8�;�&�>�}�3���0������XN�����9�u�<�;�;�}��ԜY������R�����0�&�:�u�1�2��������G	��X �����=�&���]�}�Zϐ��Ƹ�R��s��<����8�,�7�w�0����Y�����������u��;��"�)�W���ӕ��Vl�C����� �u�0�0�w�8����Y����_��Y�� ���3�7� �1�y�}��������A��~N��I����!���$�<��������_��R�����d�y�:�4�6�3����P��ƹ	��C��&���4��u�i�w�����(ە��_
�������&�0��6�2�l�[ϱ�����z��OG����x�u�'�4�2�)�Ϯ�����Z��U�����x�#�:�>�2���������c��u�����x�#�:�>�6�����:����E��[ךU���=�:�
�u��<����Ӊ��R��V�����u�x�#�:�<�<��������_��X*�����4�<��!�]�}�Z�������@"��V'�����u��!���/����Y����[	��h��1�����%��8�<��������bl�C�����4�.�&�{�~�}�S�ԜY����G/��R�����9�6�-�u�9�4�ϩ��Ȋ�R��Y�����6�9�6�u���}���Y����A��Z��]���u�u�>�4�'�8�'��� ����F�	N�����0��'�,�;�q�W���T�ƥ�F��C��ʧ�;�0�d�!�w�}�J��Y�����R�����4�!�'�u�w�c��������X ��C��U���u�x�<�u�>�)��������T��XN�O���_�u�u�u��0����
����f��DN��U���8�'�6�&�>�:����P����� �� ���u�h�d�_�w�}�������9F�N�����0�9�u�u�w�}�W���Y���F��R�����u�u�u�u�w�}�W���Y����]F��C
�����_�u�u�u��<�������F�N��U���k�:�!�'��1�0���U���F�N��X���;�u�:�9�6�W�W���Y����@�N��U���u�u�u�u�w�c����
���F�N��U���u�u�u�x�w�3�W���
����X5��G��%���,�u�u�u�$�<��������F�N��U���h�u��!���������F�N��U���<�u�7�:�2�3�W���Yӕ��G��V
�����&�3�&�!�9�`�W�������W'��E��:���0��y�u�z�4�Wϋ�
����WT��E��¾�4�_�u�u�w�����)����F�N��U���u�k�:�4�6�3�������F�N��U���u�;�u�<�9�9�F�������V�N��Uʦ�4�4�;�<�2�}�W���Y���F�������'�4��w�}�W���Y���F��N�����}�b�1�"�#�}�^���Y����r��Z!��#���1�u�u�u�w�}�J���8����|��V��Y���u�u�u�u�w�p��������RǻN��U���6�8� ��w�}�W���Y���[�X/�� ���!�y�u�u�w�}�W���Y���	��*�����
�}��8�;�.��ԜY���@'��B�����u�u�u�u�w�}�W�������^)��fG�U���u�u�u�u�w�p�W���Y����|��CF�����0��'�_�w�p�;���Ӓ��	��G��U���8�!�0��2��Ϻ�����@	��_�����u�'�u�0�2�+�Ͻ�����_ǻC����=�u�4�%�2�1�W������F��X���0��>�_�w�8��ԜY���Z ��^�����2�}�#�'�;�t����s���F�/�����:�6� ��#�<����	�ƥ�	��T�� ���9�1�4�&�%�.� ���Y����[ǻN��U���!�'�0�6�8�6����ӑ��W	��C��U���6�0�u�=�w�<�����Ƹ�^��=N��U���3�:� �%�#�$�Ǳ�����`�������!�0�_�u�w�}�W�������G0��^
�����h�:�6� ��)����B���F��[��U���u�u�:�6�"���������VF������ ��9�1�>�8����8����|��V��N���u�u�0�1�>�f�W���Y�����_N��ʱ�!�u� �%�#�}��������r��Z!��#���1�4�&�'�$�}�W����Σ�P��x�����|�!�0�_�w�}�W���8����|��^��U��:�6� ��#�f�W���Y����r��Z!��%����i�u��4�0����s���F��SN��N���u�0�1�<�l�}����	����@��N�U���4�0�!�0�1�3�Ϙ�
���F��R��3���!�4�&�0�w�5�W���	����R��U��U���!�0��8�;��Ϻ�����R��G�����!�0�1�!�w�/�Ͻ�����Tl�C��ʡ�0��u���9����ӑ��]F��RN��U����4�,�6�%�3��������W��D�����_�u�x�=�8��W�������)��a�����%�u�x�#�8�6�ϵ�����R
�IךU���=�:�
�u��.�ϸ���ƹK��_��*����u���#�(�1���Y����[	��h�����4�%�0�9�]�}�Z�������P"��X1�����<�}��6�:�(�!�������l�C�����4�6�u��4�0��������_l�x������:�o�0�#�)�W���ݢ��\��GN�����u�u�2�;�%�>����Q���F��e�����u�k�r�r�w�p�W���Y����_	��TN�U��_�u�u�:�#�0����Y�����D��H���4�&�y�u�w�}�W���Y���F�N��U���x�u�;�u�8�1��ԜY���P#��N��Kʦ�;� �%�!��q�W���Y���F�N��U���x�<�u�7�8�8����Y����_�N��U���%�0�9�y�w�}�W���Y���F�N��U���u�;�u�!��2��ԜY���P"�N��Kʡ�
�!��2�4�2����6����_��^��Y���x�<�u�&�3�1����Y�����N��H����6�8� ��1����P���F�N��U���x�u� �u�#�����Y����a��C8������;�'�!��)�8���s�ƪ�AF��T'�����;�>�4�%�2���������W	��C��U���0�4�0�u�w���������C��V��3��u�u�3�'�>�4�W���ӕ��P��B�����%��1�-�p�4�Ϲ�����Vl�N��Xǣ�:�>�0��;�-��������w��q��<���u�u�x�#�8�6�ϵ�����R
�IךU���u�x�=�:��}�%���Ӏ��@ǻN��U���=�:�
�u��}�2�������uǻN��U���=�:�
�u�;�}��������F�N����>�4�6�u��>����)����5��~ �����|�u�u�u�z�+����Ӆ��@'��B�������6�;�2�t��ԜY���|��B�����:��u�;�>�$� ���W����C"��F���ߊu�u�u�u�2�8�������F�N��Uʾ�0�0��9�j�}�G���Y����]F��C
�����u�h�r�r�w�}�W���	����^��d��U���u�u�4�0�2�}�Iϸ����F�N��U���u�u�u�u�w�}�ZϷ�Yӄ��_��=N��U���u�u��u�w�`�W���6����G ��N��U���u�u�u�u�w�p�W���Y����V��N��U���u��>�u�w�c�$�������F�N��U���u�u�u�u�w�p����
����\��=N��U���u�u��u�w�`�W�������G6��R'�����1�-�}�|�w�p�W���Y����_	��Td��U���u�u�6�u�w�}�Iϭ�����F��['�����1�-�}�|�l�}�Zϱ�ӕ��l
��^��Hʾ�0�0��9�]�}�W���T����X9��s(�����u� �%�!�6�<����s���F�A�����>�0�0��;�z�P���Y�����X��U���&�!�3�9�2�}�W���Tސ��\����U����!� ��$�}�W���Tސ��\��-��U���%�0�9�_�w�}�W�������RF������� ��%���>����Pۏ�F�N����>�4�6�u��>����5����`��Y
��\¼�_�u�u�u�"�-��������b\��Y��ʢ�'�{��:��-�_���P���F�	�����u�4�u�_�w�}�W���Y����V��[N��U��|�u�x�<�w�.�������F�d��U���u�%�'�u�6�}�}���Y���F��R��U��3�9�0�u�w�}�W���Y���F�N��U���<�u�7�:�2�3�W���Y�����N��H�����!� ��.�W���Y���F�N��X���;�u�:�9�6�W�W���Y���p
��N��Kʆ�8�9��>�w�}�W���Y���F�N��Xʼ�u�&�1�9�0�>�W���Y�����N��H����6�8� ��-�&Ǎ�����KO��B��X���;�u�!�
�8�4�}���Y���F��N��U��&�6� ��#�>�&Ǎ�����KO��G�U���:�!�&�1�;�:���Y����V��[d��Uʰ�1�2�;�'�#�}��������G��s��3���_�u�;�u�2�8����>����R��V�� ��_�u�x��$�:�W���Y����_F��E�� ���!�_�u��4�0�������F��h�����}��6�8�"���������F��T��:���u�h�&�6�"�����0���@'��B�����h�&�6� ��)����s����4��d