-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����;�!�#�1�z�}�����Ɔ�[��Z�����x�u�'�2�9�1�'�������c>��h[�@�߇x��!�o�e�}����K����KǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��t�E��Y����A��CN�����4�u�;�!�"�8��������R��Yd�U���u�<�=�&��.����s����R��Y��<���'�8�;�&��)����Y����A��^��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��)����@��:��ʳ�9�u�'�4�2�}��������@����ʳ�'�!�0�3�6�)����Y����^��E@חX���u�u�u�u��8��������TF��^��ʶ�8�:�0�u�1�<��������]�������<�<�;�_�z�}�W���Y����R
��[�����;�!�u�;��<�Ϗ�����^��E����4�u�u�;�w�}�6��T���F�N�����&��6�0�2�)����
Ӓ����C��U���6�u�:�u�"�5��������V��C��X���u�u�u�u�w�(����Y����V�� ��U���6�9�!�:�y�p�}��Y���F�������0�3�;�2�����
������D�����0�u�'�8�#�8��������[��=C�U���u�u�u�7�1�/�W����ƿ�]��_������6�:�3��1�Y�������@F��Y��ʡ�4�u�=�_�z�}�W���Y����\��^�����:�>� �u�6�}����Y����W��D�����:�u�=�u�2�2��ԑT���F�N��Uʦ�<�=�&��2�;����?����Z��tN�����!�0�6�;�%�1����Y����[��B���߇x�u�u�u�w�}��������]��_��ʷ�u�0�#�6�3�?�W���
ӫ��	��D��U���!�0�;�-�y�p�}��Y���F������6�0��;�$�3�W����Ƹ�Z��[��U���u�4�,�6�4�8�W���
����WF��R ��X���u�u�u�u�w�<��������Q��E��ʦ�;�&�!�0�'�<�Ϫ�Y����]��#��[���3�!�<�_�z�}�W���Y����r%��V�����=�1�4�9�8�}��������P��C����� �0�!�0�4�/����T���F�N�����0�<�u�'�6�8�W���ӕ��T��C-�����1�-�:��>��4�������[��z/��X���u�u�u�u�w�4�ϭ�����]����ʘ��=�&�6�:�1��������UF��DN�����4�<�;�x�w�}�W���Y�Ư�P
��d����u�u�u�u�w�6��������Z��D�����&�=�"�8�9�}��������R��R�����0�"�<�!�9�4��ԑT���F�N�����4�4�8�8�%�8�W�������R��T������!���;�9����
Ӓ��@F��X�����_�x�u�u�w�}�WϪ�Y����VF��RN�����;�u�;�u��)�>�������@F����U���4�8�8�'�2�s�2���s���F�N��U���8�;�u�;�#�8��������_��V��ʶ�'�0�%�;�$�)�W�������]��YN�����;�_�x�u�w�}�W�������w��~ ��U���u�4�4��:�/��������Z��G�����"�<�0�y� �4�ϳ�����9K�N��U���u�&�;�9�w�����0ܷ��R��RN��ʷ�u�'�!�0�w�$��������	��NN��ʰ�0�0�!�x�w�}�W���Y�ƥ���C��#���1�_�x�x�w�}�W���Y�ƿ�V��S
�����u�0�9�u�?�.����ӑ��GF��S��ʡ�u�!�'�u�2�9��������[ǶN��U���u�u�1�!�w�8����
����[��E��U���'�&�u�&�>�>��������\��V�����6�9� �4�>�3�Z���Y���F�C��U���9�7�u�:�2�?�W���Y����9K��C��U���u�u�u��6�����
����G��DN��ʻ�-�u�'�6�$�4�ϫ��ƻ�R��R��ʴ�1�0�&�!�]�p�W���Y�����E�����3�'�<�&�9�%�W���	����Z	��=C�X���u�u�u�u�w������ƭ�WF��T��<���4�0�!�0�3�)�W���Y����P	��B��U���8�!�0�%�2�4��ԑT���F�N�����&�<�2� �>�s�W���
ӂ��RF��[��ʴ�1�1�!�u�?�}��������G��U�����x�u�u�u�w�}�W������9K�N��U���u�&�6� ��)����Y����P��DN�����=�u��6�:�(�>Ͽ�ӕ��P��B�����0�u�'�_�z�}�W���Y����R
��N�����"�9�u�0�#�6�ϸ��Ƹ�VF��D�����&�<�2� �>�}�Ϫ�Ӆ��ZǶN��U���u�u�!�u�9�4��������G��Q��ʺ�!� �u�&�!�1����
����^)��~N��ʦ�6� ��!�]�p�W���Y�������U���4�u�:�%�#�9�����ƪ�\��_�����0�&�;�u�;�>�Y��s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���<�'�'�u�2�8�W������F��^��[���
�:�<�
�f�i����s�ƹ�VF��R�� ���<�
�!�{�;�f�Wϫ�ӑ��XH��P �����!�0��%�6�1�}���
�ƻ�A��\	�����:�4��6�:�)�������F��@��[����%�4�9�]�8����Y����G"��g�� ���u�&�u�2�9�/��ԜY�Ƨ�R��Y/��&���u�u�o�<�w�3����Y����VF��C��U��d�_�u�u��/��������F�N��U���9�4�n�u�w�6����4����@��T��U���<�!�2�'�l�}����Q�����R�����u�u�;�7�8�8��ԜY�Ɵ�^��t��U��<�u�!�
�8�4�L�ԜY�ƿ�[��~ �����!�o�<�u�9�4��������[��u��X���:�;�:�e�l�}�Z��W��ƹF��{�����0�3�;�0��/����8�����B �����}�d�1�"�#�}�^���T޳��W��N�����=�&��0�1�3��������~'��N��U���<�;�1�d�w�2����I���K��@����u��9��4�8�:���
����	F�������1�b�1�"�#�}�^���T޳��l�N�����!�:�3�u�w�3��������9F������=�&��9�3�}�W�������R��N�����'��4�0�w�}�W���ƹ�@��R
��;���=�&��!�z�}�������F�b\�D�ߊu�u��4��9�������	F�������1�m�1�"�#�}�^���Tӳ��
lǻN��;����6�=�&��)����Y�ƣ�GF��X���ߊu�u��-��>����6���F�N��ʠ�&�2�0�}��0����;����F��@ ��U���u�x� �f�f�W�W���
����z��[��U���;��:�0�9�8��������z��N=�����d�1�"�!�w�t�}���Y����R/��N��U���;��2�0�f�����ۍ��G��v�����x�d�1�"�#�}�^���Tӵ��WǻN��1�����u�u�m�4�W�������r��N1�����4�;�'��-�}�W�������V�C�&��d�_�u�u��<�6�������GF��X�� ���2�0�}�u�8�3���B���f_�=d��Uʦ�6� ���m�4�W������F��@ ��U���u�x�u�a�y�W�W���8����z��N��U���;�1�a�u�8�3���B���5��]װU���&�6� ��#�<����Y����Q	��R�����u��6�8�"�����Y����@��R
��Bʱ�"�!�u�|�w�p�W��W���F��T��:���6��o�:�#�.����Q����\��XN�N���x��m�f�w�}��������zF��X�����0�}�b�1� �)�W���Y���`R��d��Uʦ�6� ��!�w�}��������R��S�����|�n�u�x��e�D��Ӡ��P��T>�����!�_�4�6�>�8����Y����\ ��E��1���'�6�;�!�>�W�}���������R�����<�0�u�u�8�1����DӒ��V]ǻ�����&�0�0��>�8����
����\	��V ��Hʳ�9�0�_�u�>�3�ϭ�����G%��T*�����u�:�9�4��>����Y����G	�N�Uº�=�'�u�k�1�1���Yӕ��]��D-�����&��!�4�>�����CӤ��_��a�����u�:�;�:�g�}�J�������[�Q����u�&�2�4�w���������Z��[��Oʗ�:�0�;�0�#�/�F�������V�S�����'�u�k�3�;�8�L�ԜY����Z��RN�����u�!�<�2�]�}�Z���������CN�����&�2�4�&�6�8��������WF��C�����&�3�:�u�#�8�W�������@F����ʡ�0�u�x�u�8�)��������Z��_�����!�'�7�!�w�8�ϱ�Y����V��^�����&�u�u�<�9�1��������lǻC�����
�<�&�4�#�}�����ƿ�R
��_��:���u�;�<�;�3�6��������@��C��U���;�:�e�n�w�.����Y����P6��D�����<�o�7�:�2�3�}���������R�� ��&�2�0�}�e�9� ���Y����F��P ��U���!��8� ��}�����ލ�A��CF����!�u�|�_�w�4����
����~��B��U���;�1�m�'�6��_�������V�=N�����9�&�0�!�6���������	F��D������8�=�&��)�Z�������V�=N�����9�&�0�!�6���������Z��[T�����4�n�u�&�0�<�W���
����p��N�����;�_�u�x�?�2�(�����ƓQ��YdךU����0�!�u�?�}�����Ʈ�\��N����>�0��4�#�8�'���,����\��XךU���=�:�
�u��.����
����a��Cd��Xǣ�:�>�4�&�2�)��������G0��^
��;����6�=�&��)����5��ƹK��_��*����-��6�?�.�8���
����~��_��:���6�_�u�'�4���������p	��E��Oʰ�!�!�u�:�<���������P3��C-�����u���_�w�}�������9F�N�����0�9�u�u�w�}�W���Y���F�	N������>�u�u�w�}�W���Y���F�C�����!�
�:�<�]�}�W���+����A�N��U���u�u�u�u�w�}�Iϭ�
����@��N��U���u�u�u�u�w�}�Z����Ʈ�\
��Yd��U���&�=�&��4�8����Y���F�N��H����4�0�;�%�0���Y���F�N��U���<�u� �&�0�8�_������F��{�����0�3�;�0��/����8���F��X�����3��1�-�8�	����:���K��YN�����;�1�d�u�]�}�W���1����@��R������'�=�&��}�Iϭ�����G%��Q�����:��<���}�Z����ƹ�@��R
��Dʱ�u�u�u�&�6�>����
����@)��N��U���u�h�u��;�����4����|��N��U���u�u�x�<�w�(��������W	ǻN��U���4�!�=�&��1����Y���F�S����'��4�0�6�4�[���Y���F�N�U���u�:�9�4�]�}�W���*����c��RN��U���u�u�u�u�w�}�Iϭ�����[��N��U���u�u�u�u�w�}�Z����ƹ�@��R
��;���u�u�u�&�2�)��������G0��^
��U���u�h�u��/�����
����e��S"��Y���u�u�x�:�#�?�������F��y��8���=�&��!�w�}�W���Y���F��R�����4�0� ��;�}�W���Y���K��B�����;�1�>� �]�}�W���+����A��[��U���u�u�u�u�w�}�Iϭ�����G%��TB��U���u�u�u�u�w�}�Z����Ʈ�\
��Yd��U���&�4�6�=�$��������F�N��H����9��4�2�(�!������F�N��U���:�!�7�:�2�3�W���Yӕ��_��V�� ���u�u�u�u�w�}�W��Y����P6��D����u�u�u�u�w�}�W���TӉ����^	��¾� �_�u�&�2�)��������G0��^
��Hʦ�0�!�4��6�8��������_]ǻ�����6�=�&��#�a�W�������c��R!��9���_�u�x�u�%�<�Ϫ�Ӆ��U ��^��U���6�9�!�'�w�p��������A��s������9�_�u�z�5����Y����@�������4�0� �_�w�/��������U%��T����!�u�:�>��<����:����p��F��9�ߊu�u�0�0�>�}����s���F��X��8���;�!�;�0�j�}�4�������]��Y��U���u�;�u�;�2�8�W�������G	�=N��U���!�8�%�}�w�}�Wύ�����_�N��U���%�0�9�y�w�}�W������G��X	�����u�u� �0�;�����D�ƿ�@��C-�����u�x�u�;�w�2����s���F��_��<���u�u�k�&�6�>����6���K�^ �� ���2�0�}��:�<����
����@K��S�����|�u�u�u�$�2�������X��t�����|�u�u�u�z�2�ϭ�����T��X����_�u�x�u�>�8����
����R��V�����&�4�6�=�$������Ƹ���G�����3�'�!�0�w�p�W�������V��T�� ���<�;�1�9�.�W�W�������`��[���ߊu�0�<�_�w�}�Ϭ�
����V��=�����9�|�!�0�]�}�W���+����A��[�����i�u��&�6�)��������@4��C��6����9�,�=�0�p�W������F�D<������9�n�u�w�}��������V)��a�����4�u�h�&�6�>����6����_��R��]���9��4�0�"���������[��_�����:�e�u�u��1�'�������R
��d��Uʰ�1�<�n�u�2�9��������9F�N�����!�!�0�8�:�/�W����Ƽ�Z��EN������&�!�1�6�.����s�Ƽ�\��DF������>�_�u�2�4�}���Y����Z��P1�����4�%�0�9�~�)��ԜY���@3��E<�����%�u�h�&�$�/����B���F��e�����!��1�0�$�a�W�������V��G�����:�u� �0��.��ԜY�Ʃ�WF��d�����%�:�0�&�]�}�Z���������
��ʸ�8�'�_�u�z���������V��E�����;�u�4�6�?�.�8�������R��S�����7�u�"�u�;�>�W������2��DN��U���0�7�6� �2�)�Ϻ����K��R��ʧ�4�u�4�=�>�}� �������P��RN�����'�!�4�u�?�}��������GF��[�����;�%�!�{�w�)��������AF��
���ߊu�x�!�0�2�)�ϭ�������_�����u�0�4�<�0�)�ϻ�����z7��V��ʴ�!�'�!�0�:�0�������F�A������4�!�0��)�:����ƈ�G��Z�����x�=�:�
�w���������r��X�����'�0�u�x�!�2��������|��E�����_�u�x�=�8��W�������W'��E��<����&�4�!�6�>����Q��ƹK��_��*��� �1�!��6�����
ӕ��_��V�� ���9�1�0�4��t�W������l��e��4���0�&�;�&�2�9����
����F�A�����&�4�4� ��.��������zl�C�����4�&�4�4�"���������F��N����>�4�&�0�3�9����6����a��v
����� �_�u�4�6�8����Y����G��X��3���!�0��!��0����+���F�P�����8�%�}�u�w�}��������G1��S
�����'�h�u�'�2�}�W���Y���K�^ �����0�;�o�u�%�8�W���YӍ��G��v�����u�u�u�u�j�}�3���0����`��N��Xʼ�u�<�!�2�%�/����HӒ��F��\ךU���u��!��#�/�$���Y���F�	N�U���u�u�u�u�w�}�ZϷ�Yӏ��V�������u�:�g�o�w�W�W�������R�=N��U���4�%�0�9�w�}�W���Y���`��[�����u�u�u�u�w�}�W���Y����]F��C
�����_�u�u�u��.��������A��S����0��<�0�3�/���Y���F�C�����:�9�4�_�w�}�W�������W'��E��<���k�&�0�!�%��������J�N��U���u�;�u�:�;�<�}���Y�ƿ�C��R<�����'�&�u�k�$�<����
����e��S*�����|�u�x�u�9�}�������F�D<�����'�&��u�w�}�Iϭ�����W��D'��U���u�u�u�u�w�p�W���Y����T����G���&�}�d�u�w�}�W���
����z��[��U���u�h�u��#��!������F�N��U���u�x�<�u��2����������C��4���_�u�u�u��)�>���Y���F�S����4�;�y�u�w�}�W���Y���F�C�����<�;�1�m�%�<�(���=����]'��N��Uʦ�4�4�;�u�w�}�W���Y����w��~ ��U���u�u�u�u�w�}�W���T�ƥ�F��P ��DҔ�'�,�!�>�6�<����Y�����C�����u�u�u�u�j�}�3���4����G/�N��U���u�u�u�u�z�2�ύ�����'��V��]���!��!�_�w�}�W�������bF�N��U���k�&�4�4�2����Y���F�N��U���u� �u�<�9�9�O�������X"��V!��4���u�u�&�0�3�9����6���F������1�0�&� �~�}�W���Y���K�X�� ���2�0�}�:�e�8����H���9l�C�����0�!�0����W������l��E��'���8�9�'�4�w�<�>���Tސ��\�������!�4�6�&�2�)��������R��e�����4�6�0�4�p�4��ԜY�˺�\	��VN�����4�<�u��;���������Z��[�����6�=�&��#�<��������Z��=N��X���:�
�u��2�;�ϭ�����FǻC�����
�u��!��}�3���4����G/�d��Xǣ�:�>�4�&�4�(�>���8����z��N����>�4�&�6�"��ϭ�����F��N����>�4�&�6�"�����Y����F��C"��<����6�o�0�#�)�W���ݠ��P��D�����4�u���]�}�W�������^��d��U���>�<�&���<���Y����@��t�����x�u�;�u�8�1��ԜY�Ƽ�A��V�����u�u�4�%�2�1�W���D�Ɵ�^��t��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�p����
����F�N�����4�<�u�u�i�.��������F��[�����}��9��6�8��������_��_��\���x�u�;�u�8�1�W���Yӕ��@��C-����u��&�4�#�<�����ο�V��E�����9�,�=�2�~�}�W���Y���F�N��Uʷ�:�_�u�u�w�����Y���[�D*������!�}�|�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Tӏ����Yd��U���&�:�3��w�}�W���
����U)��N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�x�w�3�W������F��v�����u�u�h�u��>����U���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���<�u�&�2�]�}�W���8����|��N��Kʦ�6� ��!�{�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���K��B�����u�u�u�&�4�(�8��������T�� ���9�|�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�Z����ƿ�TǑN�U���4�0�!�0���4���Tސ��\��(�����&�8�9�'�6�}����Y����[	��h��'���4�!�4�6�$�8����:����V
�������!�4�6�0�6�z����s���E��\1�����4�4�<�u��1�'�������R
��s��¦�4�6�=�&��)����=������_GךU���=�:�
�u��8����
����U)��=N��X���:�
�u��#��W�������|��^��U���#�:�>�4�$�>����Y����F��fd��Xǣ�:�>�4�&�4�(�8���
����^)��fd��Xǣ�:�>�4�&�4�(�8����ƿ�P��x�����u��6�o�2�)��������A��e�����'�4�u���W�W�������PF��GN��U���u�>�<�&������D�Ƨ�Z��~ �����u�x�u�;�w�2����s���C	����U�ߊu�u�u�4�'�8����Y���`��[�����u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�ZϷ�Yӕ��ll�N�����4�4�<�u�w�c��������V)��a�����4�}��9��<����/����w��NI�����u�x�u�;�w�2����Y����a��V�����h�u��&�6�)��������@4��C��6����9�,�=�0�t�W���Y���F�C����7�:�_�u�w�}�3���0���F�	N�����0��!�}�~�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y����]F��^	��U���u�&�:�3��}�W���Gӕ��V ��B�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�z�}������ƹF������;�u�u�h�w��������F�N��U���u�u�u�u�w�}�W���Y���F�N��U���x�<�u�&�0�W�W���Y����F��CN��U��&�6� ��#�q�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F���U���;�u�u�u�$�>��������X��v������9�|�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W��Y����@��=d��X���<�0�<�0�#�8��������[��x������9�&�2�6�}�Ͻ�����@'��B�����<�{�u�=�$�>����
����9F�N��ʡ�0�6�0�3�4�8�Ͻ�����G����U���u��u�0�6�s�WϮ�����5��G�����u�7�2�;�w�}��������l��RF������>�u�=�9�}�W���
����^)��a�����4�u�h�&�4�(�8�������V
������� ��9�1�2�<�P�������\��XN�U����-��6�?�.�8�������P
��N�����<�n�u�0�3�-����
��ƹ��T�� ���9�1�i�u��>����/����w��NF������!�4�<��1�ȶ�����9��<��N�