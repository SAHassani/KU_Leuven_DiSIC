-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����0�4�{�=�]�p�6�������\��t�����x�u�'�2�9�1�'�������c>��h[�C�߇x��!�o�f�}����I��ƴl�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�u�4�}�G��:����Z�� �����9��&�'�:�3�ϝ�����G��=C�4����2�!�u�2�8����T�Ƃ�G��V����� �0�!�u�9�8����0����^��X חX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�Z�������V\�c��U���0�6�0�!�$�9��������@H��V�����0�u�<�9�$�2�ϭ�����`��=C�U���u�u�u��w�<����Wө��VF��RN����� �3�'�=�$�.����������G��U���'�1�!�0�z�}�W���Y���Q��R�����u��%�9�9���������@F�������0�1�;�u�?�}����s��ƴF�N��U����0�&�2�6�}�����ƿ�_����U���0�<�0�1�;�$����)����Z��R��8���&�<�=�_�z�}�W���Y����V��D�����<�<� �u�>�8����������G�����&�m�&�;�2�)������ƴF�N��U���%�%�9�;�w�)�����Ƹ�Z��Y��ʴ�1�!�0��#�����Y������Y���߇x�u�u�u�w�}�������KǶN��U���u�u��!�w���������]	��T��ʴ�9�!�0�%�9�4�Ϭ��ƾ�B��C�����!�_�x�u�w�}�W�������^�������;��9�,�w�<����Y����p��t�����3�0�u�=�w�<���Y���F�N�����;�4�<�u�2�2�Ͽ�
����]��e��ʢ�9�u�0�u�?�}��������@��C��U���u�u�u�9�6�}���T���F�N��U����!��,�>�8��������[��^�����=�u�4�4�5�.�_������ ��=C�U���u�u�u�>�6�<��������G��S��U���!�u�;�&�6�<����"û��R��V��ʷ�3�'�u�=�]�p�W���Y�����C��ʦ�4�4�;�z�� �W���Y����_��X��U���9� �1�!�w�3�ϩ����F�N��U����!����l�W�������l�=C�U���u�u�u��2���������@F��RN�����6�4�;�1�w�5�W���Ӊ��C��X�����4�4�7�3�2�W�Z���Y���F��DN�����&�!�0�1�#�}����Y����[��R�����0�u�;�!�2�>����Y����Z��CחX���u�u�u�u�#�}��������Q��R������!���;�9�W�������F��V�����x�_�x�u�w�}�W���
����|��V��U���4�u�'�4�w�;��������[��^ �����u�=�;�4�$�<����0ܷƴF�N��U���&�7�'�4�w�.�����ƿ�R��Y'��U���4�g�u�'�6�}����������
��ʺ�!� �&�x�w�}�W���Y�ƣ�����U���4� �3�'�w�5�Ͽ�ӂ��@��_������&�;�9�w�4�W���T���F�N�����4� ��9�3�3�W�������]��C��Uۑ�&�7�'�4�w�3��������bN��G�X�߇x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��������RB�����_�u�&�u�2�8��������lW��@���ߊu�&�u�0�2�3����������d�� ���"�'�{�>��<��������Z��X����u� �0�"�%�s����,����G��s�����_�u�&�u�8�6�'���
�ȭ�_]Ǒ{����� ���n�w�(�ϋ�0����E��G�����4�9�_�0�#�)�W�������w��s��ʼ�_�u�0�0�>�u�W�������R��B�����u�;�<�!�0�/�M���B�����C�����0�u�u�u�9�4����Ӕ��T���G��u�|�_�u�8�)�}���Y����V�N��U���9�4�n�u�w�����:�����D�����6�_�u�u�z�}��������V
�������0�{�u�u�$�4��������J+��B�����o�<�u�;�>�3�������\F��N��X��m�_�u�u�z�����Y������D�����_�u�u��1�8�$���Y�ƥ���^	����1�"�!�u�~�}�Z�W��ƹF�N�����1�!�u�:�w�5�W���
�ƨ�G��B���ߊu�u��!������Cӏ��q	��R�����'�>�4�4�%�����Y�ƨ�D��^����u��!���g��������^��E��¾�4�4�'��-�}�W�������V�C��D���_�u�u��#��&���Ɵ�T��V�����!�>�4�4�%�����Y�ƨ�D��^�U���d�{�_�u�w�p�W���	����R��Q��U���u�=�u�4�6�?����
�����C�����<�u�u� �w�2����/����AN��B�����3�0�&�x�f�9� ���Y����F�D*������o�:�!��:���8����l��y����� �3�'�u�w�}�������X"��V/��&���x�u�:�;�8�m�L��Y����l�N����� ��o�:�#�����H˧��"�������4� �3�'�w�}�W������F��V�����/�x�u�:�9�2�G���Y����^�=d��ʓ�4�!�0��#�����s����[��T��ʇ��:�u�'�4���������JF��=d�����u�;�<�;�3������ƭ�A�� �� ���u�4�2�u�i�t��������V�
�����e�n�u�!�'�}��������G	��s1�����'�4�}��:�<��������F��S�����|�:�u�:�;�<�!����Χ�R��E�����u�:�;�:�g�f�WϪ�	�ƅ�w��v��ʼ�u�'�4�}��0��������@F��@ ��U���:�u�<�;�3�e����&�Χ�R��E�����u�:�;�:�g�f�}���������C��#���1�'�u�u�8�1��������w9��=N�����9�&�4�4�"�;�������$��[��#���:�}��8�6�<�������F��@ ��U���_�u�<�;�;�.�������/��V�����n�u�&�2�6�}�3���8����	F��s��4���!�_�u�&�0�<�W�������U%��Y��U���<�;�1��.�)�FϺ�����O�
N�����&�h�u�:�"�.����Q����R'��d��Y���n�u�&�2�6�}�3���;����WF��u�����0�!�'�>�"���������W��X����n�u�&�2�6�}�%���<����VF��u�����0�!�'�>�"���������W��X����u�h�}�!�2�.�J�������l�D������4���#�5�MϜ�����e��X��;���4�4� �3�%�p�W������F��F�����u�k�3�9�2�f�WϪ�	�Ǝ�\
��C������%�
�u�$�<����Q����w��u�����d�1�"�!�w�t��������]0��C��G���1�"�!�u�~�W�W�������w��u��'���,�o��:�2�3����ۍ��^"��V,�����x�u�:�;�8�m�W��Q����A�	N�����n�_�u�x� �}�����Ư�^��D��U���u�=�u�<�2�4�Ϻ�����UF��RN�����u�:�6�0�#�}�3���6����_��N�����;�u��!��0����	����R������u�h�`�_�w�$�Ϝ�����R$��Q<�����%�
�u�&�6�/����7����G��Q����1�"�!�u�~�2�W�������V��EF�����0�:�,�<�2�8���Y����G	�UךU���;�9�&�4�6�(��������VF��u��1����3���.�4����C����G��DN��Uº�=�'�u�k�1�1����s���F��RN�����u� �3�'�?�1���Kӯ��@��[��U���!��,�<�2�9����
Ӓ����C��ʦ�0�1�1�'�$��Y�������R��\<�����'�&��0�m�(�����Π�TT��D�@��>�4�4�'��'�^Ϻ�����O���� ���2�0�}�y�8�o�B������r��^��\�ߊu�<�;�9�$�-��������W��DT�����4��6�:����������V��N�����u�|�_�u�z�+����
����R��N����>�&�2�;�]�8��ԜY����\F��[�����3�'�<�0�$�0�����Ƨ�V�������u�3�=�"�:�3�W�������R��RךU���0�<�!�:�w�5�W���Ӥ��U��!��ʡ�<�u�:�;�2�}��������G��RN�����0�&� �3�%�4����T�ƿ�^��DN��U���1�0�0�,�#�0�W���������C�����0�{�u��9�<��������F��EN������8�4�4�"�;���Y����G	�	�����0�u�u�%�8�8�Ǎ�����_�N�����;�u�u�u�>�}��������VN��Z��6���u�=�;�u�w�}�WϷ�Y����V��_��U���u�u�u�&�6�<��������ZO�
N��*���<�;�1�>�6�<��������l�N��U���&�0�1�;�5�8����DӀ��@��N��U���u�&�0�1�9�<����P���U��RUךU���u�u�9�0�w�}�W���Yӏ��@"��V'������,�<�}��)�6������F��R ךU���u�u�u�u��)�5���:�����S��1����3�� �#�4�W���=����A��M�U���u�u�u�0�3�4�L�ԜY���F�C��ʡ�0�6� �!� �1�W���Y����q��R�����=�u�0�!�#�0�W�������R
�������4�'��/�z�t�W���Y���K�V�����u�;�7�0�%�<�W�������l�N��U���&�0�1�;�5�8����Dӕ��G��Q�� ���<�u�u��1�8�$���B���F�N��'�����!�=�>�}�Jϭ�������_F��U���&�0�1�;�5�8���Y���F��Y
���ߊu�u�u�;�w�;�}���Y����C��R�����u�x��u�?�}����ӏ��A��NN��U���1�u�0�1�2�8�Ϫ��ƻ���C�U���&�4�4� �1�9����Dӕ��G��a�����}�|�>�4�6�/�$���T���R��F�����;�7�0�<�w�/��������G��^G����;�u�0�0�6�8�0�������U ��dךU����!��9�3�/���YӀ����YN�� ���!��3�0�$�l��������T��E�����u�x��%�2�8�Ϫ�Ӑ��Z��RN�����7�&�1�:�w���������R��Y�����u�&�;�u��.�W���Tސ��\��(�����6�'�g�c�8�1�3���+����Vl�N����>�4�&�u��)�5���+�Υ�9F�C�����
�u��%�;�3�3��� ����@2��R��%���9�;��9�.�4������ƹF������u��&�4�6�(�����Υ�9F�*�����<�0�u�;�>�$� ���W����G"��d��@ܗ�:�u���]�}�W�������R�=N��U���u�4�%�0�;�}�W���Y���F�S�&���9��>�u�w�}�W���Y���F���U���
�:�<�_�w�}�W���)����Z��R��8���&�=�0�u�i�.��������_��^ ��0���!�u�x�u�9�}���������Y��E���u�u�u�&�w�}�W���Y���F�N��U��u��!��1��_���Y���F�N��Xʼ�u�7�:�0�9�}�W���Yӕ��F�N��U���u�u�u�u�w�`�W�������U4��[��\��u�u�u�u�z�2�ϼ�����9l�N�U���<�<�<�9�-�}��������V��NI�����u�:�;�0�w�8����Y����@��Cd��U���u��4��6�����
����]��b�����4��1�0�$�<�W���Y������RN�����u�u�x�u��.�Ͽ�
����l�N�����0�0�1�1�%�.�_���E�ƿ�V�������4� �3�1�;�u�^�ԶY���F��RN�����;�u�0�4�w�3��������JF��[�����&�_�u�u�z�
�W���������V��:���#�9�1�!�6�}�������@F��[��ʢ�!�u�0�%�4�}����Y���@"��V,�����9�{�u�u�'�2����*����V%��d��Uʷ�2�;�u�u�w�4�W�������W��d�����>�u�=�;�w�}�W���
����q��e
�����0�<�u�h�$�<��������J6��RF��]���!��3���$��������T�
�����e�u�u��#�����=����]ǻN��U���u�3�_�u�w�3�W�������9F������3��!�4�>�u�^��Y����R$��Q<�����%�}�|�&�6�<��������Z��^G�����n�u�0�1�0�3����Y����R��V��4���,�_�u�x�w�.��������Z�������u�3�!�0��)�W������F��V�����<��,�e�w�`��������_��=N��1����,�}�|�k�}�3���0����F��V�����e�u�h�&�6�<���s���"��D�����u�=�u�4�6�����
����_��R�����=�u�0�:�>�.�}�������@��V�����4�<�o�u�1�/�Ϸ�Y����w��u�����x�d�1�"�#�}�W�������9F�������9�1�'��t�K�������@F������3��!�4�>�u�Z���B����]��R ������;�4�&��<��������W]ǑN�U���4�0�!�0��)�W�������V��Nd��X���0�<�&�4�#�<�Ͽ�?����w��V�����,�6�;�<�"�8�W�������^����U���!�u�:�;�2�}����s�����_N�����u�=�u�0�3�-����ӂ��A��Y�����,�!�8�u�2�<����Y����R$��Q<������<�_�u�z�*�ϩ�Y����	��R�����3�'�!�u�?�}����Y����R��RN��U���'�1�<�u�3�/����WӲ����Cd��X���4�%�0�<�w�)�����Ƹ�VF��P��ʴ�1�0�&�4�3�.�W���Y����	��[����;�<�2�:�]�}�Zϵ�����J5��RG�!���'�4�u�;�w�/��������A��E�����'�0�u�3�2�}�%���Ӈ��V��d��X���=�u�0�1�'�4�����ƾ�@��C�����n��!�'� �4����
����V��M�����0�u�;�u�6�)��ԜY����c��[��1���,�<� ��0�)�����Ƹ�VF��E�����u�0� �&�w�4�Ͽ�
��������ʴ�1�0�&�%�>�)����T�ƻ�_
��G
��ʡ�u�y�3�;�;�$�W���Ӆ��_��V��ʡ�0�4�&�'�>�3�����ƾ�R��R�����;�u�x�u��)�5���+�������� ���;��!��#�}�Ϩ����F��Y*�����3�'�o�u�1�/�Ϸ�YӍ��^"��V,�����x�u�:�;�8�m�W�������9F�C�����
�u�'�6��>��������"��V'�����_�u�u�x�?�2�(���0����^��`�����;�0�u�4�$�W�W���T����X9��\*�����'��/�u��)�6�����ƹF������u��!��#�/�$���Y����R'��d�����u�x�=�:��}�%�������V'��E��U���&�!�u�u�z�+����ӕ��R��V
�����&�;�&�0�2�W�W���T����X9��D;�����0�1�1�'�$�}�"�������W'��E��]���u�u�x�#�8�6�ϭ�����W��D'�����1�1�'�&��8�W���Tސ��\��������9�1�&�6�<���������N��Xǣ�:�>�4�&�6�<����=����A��^GךU���x�=�:�
�w�����(ӕ��G��N?��\���u�x�#�:�<�<����������C�����~�|�u�u�z�+����ӕ��G��C?��1����,�}�~�~�}�W������l��e��4���0�&� �u�'�3�W���=����]"��V����!�u�:�>��<����=����V��NN��!���u�u�u�2�9�/�ϳ�	��ƹF�N��<���0�0�!�'�3��������U��RB��U���u�u�x�<�w�?�������G��=N��U���u��!���$����Y���F�	N�����'��/�y�w�p��������V��V ��U���:�g�o�u�]�}�W���Y����R)��v�����u�u�u�u�i�6��������VO�C�����;�0�0�u�6�:�W������F��N��Uʥ�'�u�4�u�]�}�W���Y����_��\N��U���u�u�k��:�1�4���Y���F�N��U���<�u�&�1�;�:����Y�����D������1�0�&�j�}�%������F�N��U���u�x�u�;�w�2����s���F�D"�����1�1�'�&��}�Iϭ�����F�N��U���u�u�u�x�>�}������ƹF�N�� ���!��4��3�8���Y����R��R�����&�}�|�u�z�}��������]l�N��Uʦ�0�1�1�'�$��W���Y����a��v
�����;�y�u�u�w�}�ZϷ�Yӓ��Z��SF��ع�&�d�`�g�x�6����Y�����C��#���1�u�u�u�j�}�3���0����Z��NF��Y���u�x�u�;�w�2����/����AN��V������/�_�u�w�}�W�������F�N��U���k�&�4�4�%����Y���F�C�����2�0�d��/��������z��N=��U���u�u�&�4�6�3�W���Y���F������,�}�|�u�w�}�W���Y����]F��^	�����'�4�
�}��)�>��� ��ƹF�N��1����!�u�u�w�}�W��Y����R'��~F��D���u�u�u�u�z�}��������^��E��¾�4�4� ��.�W�W���Y�ƿ�R��B��U���u�u�u�k�$�<����(ۏ�J�N��U���x�:�!��0�8�Fן�������C������u�u�u�w�.��������@)��N��H���%�;�n�u�w�}�W���Y���F���U���<�;�1�9�0�1���L�����=N�����0�0�4�0��3��������@]ǑN�U���<�;�!�0�8�)����Yӕ��G��C8�����h�&�4�4�"�;��������F��Y*�����g�o�u�3�%�4����7����G��Q�����d�u�:�;�8�m��������F�p����� �d�o�u�w�;�ϴ��Ƨ�R��E�����u�u�:�;�8�m��������F�N����� ��<�?�w�`���������F��N���u�u�&�4�6�(�&Ƿ������C�����~�|�?�n�w�}��������R��p����� �d�n�u�2�9��������t��V�� ���n�0�1���W