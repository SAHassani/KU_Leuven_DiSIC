-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:� �<�{�?�W�Zϟ�����,��YN�����4�u�;�u�8�8�4�����ƴF��^	�����'�?�6�o���(��L���"��RT��Bʟ�9�u�e�d�z�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��C�����e�d��%�%�:�ϐ�����_F��D�����&��'�:�6�4���Y����a��C�����#�1�x�u�6�4����0����F��C�����;�9��3�%�<����T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x�u� �%�$�g�W���
Ӌ��F
��T�����:�0�%�:�2�.��������\��_�����<�;�9�x�w�}�W���Y�ƥ�G��X�����x�_�x�u�w�}�W���-����^	��[�����&�4�;�"�4�1��������E����ʦ�!�'��9��W�Z���Y���F��D�����u�!�"�9�w�<�����Ƨ�E��[��3���:�u�:�3�>�4��������9K�N��U���u�:�3�:�w�����Ӈ����C��ʡ�0�u�<�=�#�8��������W��
��ʼ�u�=�_�x�w�}�W���Yӕ��U��R	�����{�x�_�x�w�}�W���YӲ����T����� �<�u�<�;�<�Ͽ�Ӊ��G��Z�����u� �%�!�w�2�Z���Y���F�D/�� �����!�u�%�<�Ϫ�ӕ��P��B��$ʺ�!� �u�=�#�4�W������F�N��U���=�;�&�6�"������ƭ�@��D@��;���1�!�u�&�$�4��������G��D�����u�u�u�u�w�}��������Q��D�����u��!���1�ϩ��ƺ�_��S��U���u�,�9�&�z�}�W���Y���_��EN��U���!���%���}��T���F�N�����4�4�<��w�3�����ƥ���E��ʻ�"�1�!�u�8�?�W�������]��C�����'�0�_�x�z�}�W���Y���u	��\=������'�,�9�w�}�[ϭ�����R��S�����&�!�;�6�9�<����ӏ��V��=C�U���u�u�u�:�1�8�W���Ӓ��Z��E�����<�&�u�4�'�8�W�������[�������'�n��<�w�.�Z���Y���F�Y�����0�4�&�u�2�}����������P�����3�>�4�%�2���������[�����߇x�u�u�u�w�}����ӂ��RF��YN��U���=�1�!�u�?�}�������V����ʼ�u�&�;�!�.�)�����ƪ�Al�N��U���u�u�=�u�"�/��������R��Y@�����u��!��6�����
����V���� ���4�0�w�e�{��F�ԑT���F�N�����d�w�_�x�w�}�W���Y���F�;��U���u�0�0�!�3�)�Y�������GF��X�����4�!�#�9�3�9���T���F�N��U���u�u�<�6�"�4�ϰ�ӂ��RF��R ��1�����9�1�6�.����W���F�N��U���e�u�k� �2�)�ϭ�����]��D�����u��0�0�#�m�����Ơ�@��V��U���4�_�x�u�w�}�W���Y���F��Y�����u�0�u�4�6�*����=����]0��^
�����!�|�_�x�w�}�W���Y���F�;��U���u�=�'�u�2�8�Ϻ���ƴF�N��U���u�d�u�k��4�W���������^
�����!�_�x�x�w�}�W���Y�ƛ�V��R�����<�u� �=�3�)�W���Y������C�����u�<�0�4�9�*��������\ǶN��U���u�u�&�4�#�}��������GF��C�����=�u�4�!�3�)�W���ӑ��_F�������u�:�!�0���}��Y���F������3�9�:�<�0�6��������p��RN�����{�x�_�x�w�}�W���YӲ��@F��P ��U���!�8�u�9�0�8�W���
����e��S'�����x�u�u�u�w�}�W���Y����GF��P ��ʴ�0�0�%�6�2�}�϶��ƨ�U ��R �����9�;�u�0�6�.�}��Y���F�:��U���9�"�;�u�6�<����
ӂ��P��RN��ʧ�$�<�0�0�#�;�ϻ��ƿ�T��d����u�u�u�u�w��W�������P��R�����3��9��'�����Y����R
��[��U���u�:�3�<�>�3���Y���F�N�����&�!�'��;��W�������2��DN�����!�0�6�'�2�-����ӂ��RF��EN�����u�u�u�u�w�}��������]F��R
�����0�6�u�=�w��W�������_	��DN�����u�3�0�_�z�}�W���Y����`��C-�����4�&�'�&�w�)����
����J��DN��U��� �0�:�!�#�8����ӂ��Rl�N��U���u�u�0�:�.�/��������@F��B��U���9�u�:�'�6�}����������VN�����0�:�,�_�z�p�W���Y���F��V�����<�u�;�u��)�%���8����@��Q��<���=� �1�x�w�}�W���Y�ƫ�GF����ʠ�<�u�u�>�6�<����=����F��T��U���0�u��4�#�<����s��ƴF�N��U����u�4�0�w�*�W�������\F��^�����!�0�u�0�3�9��������[��e"������8�'�0�{�p�W���Y���F�������=�u��0�1�<��������JF��V�����0�z�u� �#�5��������W��=C�U���u�u�u�c�4�2���� ������R��&���!�4�6�;�6�.��������]��[��U���9�u�3�0�]�p�W���Y�����C�����;�_�x�x�w�}�W���Y�ƿ�G��t��:���u��4�0�"�q��������R
��N�����0�1�1�'�$�����6����]ǶN��U���u�u�&�4�6�(�'���0ܷ��A��[�����<�0�u�0�$�2�ϱ�Y����P	��R�����2�<�%�!�z�}�W���Y���@��V�����u�=� �1�5�}�����Ƹ�VF��O�����&�<�2� �>�s�W���
�ƿ�T��Dd�U���u�u�u�u�%�}�����Ʈ�-��R�����4�!�'�6�4�8�W�������]��X�����6� � �4�>�3���� ���F�N��Uʺ�u�=�u��w�3��������r%��^�����0�&�=�&�w�2�W�������P��T��U���9�&�4�1�z�}�W���Y���R��Z�����9�u�=�u�%�9����W���K�N��U���u��6�;�#�3�Ϻ�����]��@��ʶ�0�3�6�0�#�}����
����JF��^חX���u�u�u�u�>�.����W�ƚ�_��A�����4�2�u�'�:�m����7����\��D�� ���&�x�d�_�z�}�W���Y����~��Y�����<�u�9�:�"�8�W�������_����U���'�6�u�0�3�<����
Ӏ��9K�N��U���u�!�0���.�W���Ӓ����E��U���4�<�u� �#�-��������Z��T�����;�<�2�x�w�}�W���Y�Ư�V ��T�����_�x�u�u�w�}�Wϊ�Ӏ��_F��G�����0�4�u�=�8�:�W���
Ӌ��F
��^��%��� �<��6�:�8��ԑT���F�N�����&�_�x�u�w�}�W�������f��c�����4�u�h�>�8�;�4���)����V
��E��8���<�0�0�4�w�}�'���,����P��s���߇x�u�u�u�w�}�W���Y���F�N��U���h�d�u�u��8��������\�CחX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�1���� ӏ��VJ��X�����&�u�0�0�$�9��������H��[UךU���u�0�0�;�:�/����݇��l�B�����{�>�� �>�4����
�ȭ�_]ǻ��U���>��2�&�y�1�L�������\��g������!�'�{�;�f�}��
����V�������!�
�3�_�>�/��������p	��{�����'�'�u����}���Y����z+��T�����!�{��n�z�}��������G��D�����_�0�!�!�w�/��������A	��Y���ߊu�0�0�<��}�Wϵ�����@6��t����<�u�;�0�2�}����Y�Ƹ�T�
N����u��0�6�8�6��������]F��C��ʧ�;�0�g�!�w�}�J��s���X+��~ �����u�u�;�0�2�}�J��B����\��=N��U���%�0�9�u�w�3��������lǻN��&���!�4�6�;�m�4�W�������9F������;�u�u�;�"�.����Q����@��Y	��U���u�:�;�:�g�f�Z���K����9F������4�6� �u�w�(�W�������9F������ �u�u� �w�3����ۍ��R��R �����d�1�"�!�w�t�W��,���9l�N�U���u�:�9�"�9�}�����ƿ�\�������,�1�`�6�4�8�W���Ӕ��C��=N��U���!�u��4�#�<����Y����w��~ �����o�<�u�:�;�<�L���Yӕ��G��V
�����&�3�&�!�9�g��������V�
�����e�n�x�u�e�o�W���T�ƿ�R��Y>�����u�=� �1�4�3����������VN��ʶ�:�>�u�u�z�}����
Ӈ��V��d�����6�;�4�&�%�.�}���Y����R/��^��U���;�&�2�0��j��������F�=�[�ߊu�u��!������Cӏ��@��R
��Bʱ�"�!�u�|�w�p�$��H���F��V�� ���9�1�o�:�#�?�������F��V�����1�'�&��1�8�8���CӉ����^	����1�"�!�u�~�}�Zϋ�W���F��V�� ���o�:�!�&�0�8�_������\F��N�U��{�_�u�u��)�8���Y�ƣ�GF��P ��]��1�"�!�u�~�}�Zύ�A��ƓF�D/�� ����o�<�u�>�3���Y����G	�U��X���a�{�_�u�w���������Z��^	����u�:�;�:�g�f�W��*���9l�N�U���6�8� ��;�r�W�������]
��U�����6�0�u�:�$�>����0ܷƹF�N��U���,�6�8�u�8�0�Ϛ�)�މ�R��V�����;�0�u�:�0�}�Ͽ�Y���F��^	������a��6�:�2����s���@'��B������o�:�!�$�:����Nӂ��]��G�U����m�l�u�w�.����6����_7���U���;�1�a�u�8�3���B���5��WװU���&�6� ��#�<����Y����Q	��R�����u��6�8�"��Mϱ�ӕ��]��Y�����:�e�n�u�z��O��Y����r��Z!��$��:�!�&�2�2�u�@Ϻ�����O�N�U��{�_�;�u�%�>�>�������P3��CUװ���<�0�!�'�w�	�W���?����z��E�����<�u�&�_�w�2�����Ɵ�%��rd��Uʥ�'�u�_�u�w�}����Y����G��X	��U��r�r�_�u�w�}�W���ӕ��l
��^��H��r�_�u�u�w�8�MϷ�Y����_	��TN�U��n�u�u�u�6�g��������T��A�����u�:�;�:�g�f�W���Yӗ�	����*���<�n�u�u�w�,�F������G��X	��\�ߊu�;�u�:�'�3���s�ƿ�T�������1�1�'�&�w�g��������F��@ ��U���u�u�u�u�w�}�W���Y���F�T��]���0�&�h�u�g�t�}���������[<�����'�&���w�}��������E��X��U���;�:�e�n�w�p�W���Y����R��R��]���<�&�u�4�w�}�����ƺ�_��X��D���0�=�#�u�8�0������ƹK�@�����0�0�u�:�9�}�Ϫ� Ӓ��R��D��U���=�'�4�1�2�.�}���TӲ����^��U���u�1�'�&�w�.�Ϸ�Y����A��R
��ʡ�0�3�9�:�>�:��������9F�N��¾�<�!�'�4�6�8����Y����A��T�����u�u�4�}��)�%���8����@��Q��<���x�d�u�x�w�<�W�������W'��E��:���0��u�4�>�}���s���+��������9�0��#��������� ��\��:���g�u�:�u�/��Y���T�Ɓ�KF��E�����1�0�&�3�%�o�W�������T�\��U���u�u�u�d�w�p�W���Y����a��v
�����3�'�f�u��4�W��J���M�C��U���d�_�u�<�9�1��������\��T�����:�<�
�0�#�/�F�������V�=N�����9�&�4�4�"�����Cӕ��l
��^�����'�d�u�:�9�2�G��Yӕ��]��D*������!�u�u�>�3���Y����G	�N�Uº�=�'�u�k�p�z�L���
����_F��V�����!�u�u�<�9�9�F�������V�S�����'�u�k�r�p�f�}�������]��z�����0�4�u�u�w�}�W�������	[�d�����!�;�u��8���������_��N�����'�o�u��2�>��������K�d�����!�;�u��8���������_��N�����'�o�u�u��8��������w��Nd��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u��>��������F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u��:� �>���������9l�D������4�!�4�4�8����CӤ��_��a������:� �<��)�������F��@ ��U���u�u�u�u�w�}�W���Y���F�T��]���0�&�h�u�6�.�^�ԜY����R
��g�����4�u�u�u�m�����ۍ��V��X�����'�x�d�1� �)�W���Y���F�N��U���u�u�u�u�w�`�_������F��C����u�e�|�n�w�.����Y����R0��^
�����u�u�:�9�6�����Q����A��T�����u�u�u�:�9�2�G�ԜY���F�N��U���u�u�u�u�m�}������� ��D����<�;�9�&�6�<��������w��NN��U���<�;�1��%�$�ǵ�����\��V�����d�1�"�!�w�t�W���Y���F�N��U���u�u�u�h��)����D����G��DN��U��|�n�u�&�0�<�W�������_��T�����1�m�'�4��u�8�������u��X��U���:�;�:�e�]�}�W���Y���F�N��U���u�o�u�:�?�/�W���Q����A�	N��R���_�u�<�;�;�.����=����F��d�����'�,�!�<�+��������G	��N����!�u�|�u�w�}�W���Y���F�N��U���h�}�!�0�$�`�WǱ�����X�I��N�ߊu�x��6�w�/��������Z��G�����<�3�'�;�w�2��������F��SN�����:�3�<�<�9�W�W������\��R�����4�4�u� �?�4�W���Y����A��QN��U���u�<�!�'�w�$����ӇƹK�S�����!�>�<�!�%�<�����ƣ���_N�����&�;� �<�w�8����Ӄ��[F��R�����!�u�x�u�>�5����������V��ʡ�0��!�{�w�>�����Ƨ�Z
��E*�����4�u�u�;�2�8�W������p
��\(������>�4��$�<���s�����[<�����'�&�u�&�4�1�����ƪ�\��@�����&�u�:�3�0�/�W���Y����^�������x�u�0�;�2�}�����Ƣ�]K��Y�����4�!�"�u�6�}��������[��X �����%�'�u�'�:�)����T�ơ�K��ZN�����'�&�{�u�z�}��������R��E�����&�u�;�9�$�.� ����ƭ�@	��V�����u�=�u�4�>�(�}���Tӕ��G��V
�����&�3�&�!�]�}�Zϳ�ە��G��V
�����&�3�&�!�w�}����=����V��S
�����3�0��|�z�6��������w��Nd��X���'�u�x�u�6�u�3���+����W��D�����|�h�>�#�%�1��������F��OF�����0�1�1�'�$�����0���WǻC����4�0�1�1�%�.�8������X)��E�����6�:�u�u�]�}����ӕ��G��V
�����&�3�&�!�m�(�����Π�TT��D����'�9�6��4�2�W���Pӂ��]��GךU���u�u�u�u�w�}�W���Y���F�N�Uº�=�'�u�k�p�z�L�ԜY����R
��t�����o�&�2�0��o��������lǻC�9���!�!�0�8�/�;�±�Ӊ��G��D�����!�4�u�'�w�2����ӄ��F�������_�u�x�%�6�8�W�������G�������0�!�'�u�6�<����
���R��^��ʸ�-�3�;� �m�.����B����G��U��U���
�4�:�!�8�}�$�������W��DN����4�u�&�w�u�W�W�������VF��O1�����u�3�&�4�6�<���������Y�����l�n�_�u�z�5��������AǻC�����
�<�0�1�]�8��ԶY���p��C�����=�&�u�;�w�<�Ϻ�����V��C�����x��0�:�#�(�ϱ�Y������[N��U���!�!�u�=�w�8�Ϯ�����Z��B ��[���%�:�0�&��0�������Q��Yd��Uʼ�u�<�<�2�2�:�_���	����XO��_��U���u�&�=�&��1����Y���@6��D�����&�=�&��;�$����T�ƨ�D��^��Sʦ�=�&��n�w�}�Wϭ�����R��Q��1���,�i�u�&�6�<��������w��NF�����0�1�3�&�#�8���������Y��E���u��!��6�����
����V��d��U���&�4�4��;�$�K���
����z"��V��1����0�4�r�>�5�FϺ�����O�������%��_�w�}�W�������_��S�����4��9�,�$�<��������Z��N�����u�|�s�&�6�<������ƹF��Y
���ߊu�;�u�'�4�.�L�ԜY����R4��S/������3�0��#�a�Wϭ�����R��Q��1���,�>�#�'�;�>�1������O��N����� ��i�u��)�>����Χ�E��[��3���:�u�u�|�]�}�3���6����[��s��$���4�}��0�4�2�������W�=N��%���0� �u�h�$�5��������|��T�����!�'�x�d�l�W�W��-����R��B�����u��!��6�����
����V����G���7�'�u�<�"�<����Y����[��^�����'�0�_�u�z�.����
����A��[��*���_�u�&�0�#�.��������W��D!�����;�i�u�_�w�}�����Ŀ�R��R�����&��3�0��}�Ϸ�����F����U���0�4�0�4�w�3����Y����R��R��]���4�0�u�=�9�n�U���
����Z��R���ߊu�x�&�;�?�.�Ϫ�����G��YdךU����0�!�u�?�}����Y����F
��^�����,�'�2�&�2�.�W��Y����]��Z�����#�9�0�:�w�5�Ϻ�����@F��Y��ʡ�0���!�w�8����Y������B�����_�u�'�6�$�u��������9F��R	�����u�3�'�&�9�����*����V%��N���ߊu�u�u��6�)��������[�D=�����9��9�,�$�)��������R��^	��Dʱ�"�!�u�|�q�.����:����]]ǻN�����3�_�u�;�w�/����B���F�������1�4�0�#�;�8��������V
�������&� �0�u�8�.��������V��g�����;� �<�_�w�p��������\�c��U���4�u�4�6�2�}��������]��_��U���4�&�_�u��<��������[�D=�����9��9�,�<�+��������G	��N�N�ߊu�x��0�#�}��������R
��
�����0�<�!�'�]�}����
�Ο�^��t�����0�<�_�u�w�;��������T��V�����|�!�0�_�w�}�W�������Z��[��I����!��9�3�8����=����R
��s��ͽ�2�x�u�:�9�2�G���Y����R/��V��N���u�0�1�<�l�}����	����@��N�U���<�!�'�0�>�)�W����ƣ���DN�����6�4�;�"�;�}�ϭ��Ƹ��� ��ʥ�:�0�&�;�w�3��ԜY����R)��a����u��!��;�9����Q����A��T�����u�u�|�_�w�p�W�������[��s��'����1�0�&�1�.�ϝ�����9F�N�����&� �0�u�8�.����Y����[F��C�����!�0�1�!�w�5��������V��V�����u�:�!�0���}���T����|3��r<��!��� �t�&�4�6�8��������U ��CN�����u�=�;�0�>�0��������U��
�����1�;�_�u�z�)�Ϙ�>�ƥ�R��U�� ���&�!�'��;��W�������\F��[�����&�4�&�3�;�8����
����R
ǻC����>�6�6�0�w�;����+������D�����{�u�%�:�2�.�$�������l�U�����u�<�u�<�>�:����Q����_��\G�����u�u�x�u�2�(�ύ�5�Ƹ���E�����4�4�u��$�<�ϫ�����U	��C�����:�&�u�<�$�}�Ͻ�Ӕ��@ǻN��Xʡ�0�&�8�u�6�<���� Ӓ��VF��C��6����u�&�0�#�}�Ϯ�����TF����U���=�u�1�'�$�s�W���T�Ɵ�P	��N��U���u�,�9�&� �8�ϭ�����R
��YN��U���u�0�"�;�w�2����Y����]�������_�u�u�x�>�}�������g	��XN�����0�6�;�&�:�1�W�������	����ʡ�0�'�4�u�3�/�������K�G��U���0�u�4�%�2�<�ϵ��Ƹ�VF��Z�����&�{�u�u�z�}����8�Ʃ�C��DN�����9�6��6�8�}��������[��[
��ʺ�u�=�8�:�w�5�W����ƿ�G��t��<�ߊu�u�x�4�$�/�ÿ�Ӎ��V��X�����'�d�6�;�2�(����
����V��Q��U���u�<�&�u�9�s�W���T�Ƙ�V��X�����9�u�=�u�6�<�����ƥ���R��U���'�1�<�u�?�}�%������Z�������_�u�u�x�#�8�:�������F��^�����1�<�u�1�%�.�W�������W'��E��:���0��u�u��8�4�������\�_ךU���x��u�=�w�)�������Z ��R�����0�u�'�u�2�3�W�������\F��RN��9ʴ�u�=�u�4�2�)���Y���F��V�����1�'�&��1�8�>�������R��S�����!�!�u�6�8�3�W���Y����@��[�����u�'�_�u�w�p�����Ƹ�VF��Z��U���{��0�;�:�8�W���
����V�G�����u�&�>�4�'�8�'��� ����F��=N��U����0�3�'�#�8����Ӓ��+����ʠ�0�<�u�!�%�9��ԜY�����C�����1�0�&�3�$�)��������p
��\(�����x�d�x�}��0��������_�_�����u�x�:�u��)�%���8����@��Q��<���u��0�6�8�6��������`��[�����6�0�_�u�w�p� ���Y�Ƣ�DF��[�����;�&�4�!�w�8����Y����V��C�����!�0�0�0�#�)�ϓ�:ӑ��_F��R@ךU���x��!�u�?�}����Y����V��^�����9�0�!�1�#�}�������F�^��&���!�4�6�0�6�u�4�������c��s����u�=�;�u�w�}�W��Y������V�����"�<�<�2�9�*����Y����]��D�����0�<�u�!�%�9��������@F��=N��U���u�x��0�;�.�W�������G��z/�����u�&�u�&�$�2����ӕ��G��V
�����&�3�&�!�9�}�W���Y���g��R��ʡ�0�3�'�!�2�8��������r%��O�����&�&�:�0�w�3������ƹF�N��Xʦ�4�4�0�1�3�/��������]F�\!�����6��6�:�w�}�Y���Y�����Y�����4�;�4�<�w�5����Y���F��s��'����1�0�&�1�.���Y����R4��S/������3�0��w�}�8�������u��X��U��_�u�u�u�w�p� ���Y����G�������u�4�4�<�#�}����+�ƣ�VF��T�����'�u�0�&�6�)�������G��Y���ߊu�u�u�u�z�.����Y������@�����!�u�=�u��}�W���Y����V��Q��U���'�4�u�=�w�4��������Gl�N��U���u�:�u�=�w��Y���Y���K�D*�����4�<�u�0�$�)�W���
Ӄ��Z��X �����0�7�3�'�w�����)����7�D��ʶ�;�u�u�u�w�p�W���Ӏ����=��U���!�{��0�w�8����Y����U��CN�����!�3�'�!�2��4���*����V��E-�����u�|�u�u�w�}�Z�������@F��RN��ʬ�!�<�u�=�w��[Ϫ�Ӵ��WF��S��ʻ�0�&�!�u�#�/�}���Y���V
��=N��U���u�u��!��<�6�������U��R�����4�0�1�1�%�.�8�������F��A������6�:�u�w�����
����J��d��U���u�0�1�<�l�W�W���Tӯ��RF��@N�����4�<�;�<�w�2�W���������DN�����u�=�u��w�%����Y����]��
�����u�x�u�9�:�3�W�������a*�~��ʥ�&�u�0�u�6�<����Y����`4��C��U���9�y�!�0��1� ���s���K��V�����u�3�!�0�9�8��������]�^��ʴ�0�;�!�%�$�4�ϰ�ӂ��RJ��RN�����!�0�u�u�z�}����
�Ƹ���SN��ʻ�-�u�9�8�9�}�Ϫ�ӵ��l�N�U���0�"�u�0�'�.��������W��D!�����4�u�u�=�9�)�����ƿ�^��^�����:�!�;�"�4�1��������F�C�����u�<�>�1�8�s�#���Y����@��[N�����0�1�;�!�$�<��������V��Q��ʡ�u�0�'�;�>�:�W���T�ƪ�V��N��[����&�!�_�w�}�W����Ƣ�GF��V�����<�u�;�u��)�%���8����@��Q��U��e�!�0�_�w�}�W���Y����R4��S/������3�0�u�j�.��������W��D!�����x�d�_�u�w�}������ƹF�C�3���&�u�=�u��}����
�Ư�_��V��ʷ�u�1�<�2�#�8�����ƨ�_��V �����;�_�u�u�w�p����Y����G	����ߊu�u�u��;�8��������[�\(�����4�4�0�4�]�}�W���Y���F�N��U���~�'�&�/����������A��x������9�0�1�3�/��������]ǻN�����3�_�u�0�3�-����
��ƹK�t�����=�u�4�4�:�0����+�ƾ�R��S
���ߊu��9�0�3�9����*���F��S1�����#�6�:�}��1��������@O��=N��Xʒ�;�'�!�u�?�}�&Ϻ��ơ�^	��R�U���&�u�'�u�:�1�����ƻ�G��e"�����4�0�'�&�"�>��ԜY����a*��=N�����u�;�e�!�w�j��������F�C�������f��w��4���0���K��_��*���9�u�4�%�2�1�}���Y�˺�\	��VN��Uʦ�4�4�;�<�2�u�^���Y����[	��h�����:�&�1�:�>�u�3���/����w��NF�����;��0�4�w�}�3���/����w��NN�D���u�u�x�#�8�6�Ͽ�Yӕ��_4��S/�������u�u�z�+����ӗ���C�����7�}�|�u�w�p�������� W��G��U�����f��m��;��<���F��X�����}�u�u�u�w�>���Y����_��\B��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F��=N��U���u�u�u�k�$�<��������zO�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�ZϷ�s���F�T��H���:�&�1�:�>�u�3���/����w��NF�����;��0�4�w�}�3���/����w��NN�D���u�x�u�;�w�}�W������F��E�����1�0�&��{�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�C��ߊu�u�u�u�w�}�Iϭ�����G%��U'��\���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y����Fl�N��Uʤ�d�h�u�%�9�f�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�z�}��ԜY���E��\N��9���u���e��W���Tސ��\����U���%�0�9�_�w�}�Z�������WF�D*�����<�0�}�|�w�}�Z¨������������:�<�}��#���������X"��V'��$���4�u�u��#���������F��d��U���#�:�>�4�6�}����+����W��D��#���u�x�#�:�<�<����
����|��X��]���u�u�x�#�8�6�ϯ�HӉ��]l�N��9���o���d��W���YӖ��GF��GN��U���u�u�6�>�j�}��������F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W��Y��ƹF�N��U���k�&�4�4�9�4����P���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�x�>�W�W���Y�Ư�F������:�<�}��#���������X"��V'��$���4�u�u��#���������F��B��X���;�u�u�u�w�<�W��Y����a��v
������y�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F��=N��U���u�u�u�k�$�<����:����/�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�Zϱ�s���F�F]�H���%�;�n�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�x�u� �w�8�Ϲ�����VF��Y=���ߠu�x�u�<�2�4�Ϫ�ӵ��	��G��U���<�%�:�0�#�0��ԜY����V��d�����>�_�u�0�>�W�W���Ӕ��Z��R
��]���%�0�9�|�#�8�}���Y�ƿ�R��R�����h�&�2�0����������zO��N��Uʦ�4�4�0��#�}�Jϭ�����@"��V!��6����n�u�u�2�9���YӃ����T��N�ߊu�x��0�#�}��������P��CN�����4�<�;�7�8�6�W������l��E��<���'��0�3�6�>�W������l��e�����4�6�&�!�%�����s���E��\1�����3��!�&�8�;�8���K�ƨ�D��\��Uʓ�4�!�;�0�'�2��������V��C������4�!�;�2�-����:����4��d��Uʲ�;�'�6�8�'�u�W���YӍ��V��X�����'�h�u��2�>��������F�N��Uʼ�!�2�'�'�9�8�EϪ�Y����UǻN��U���6�;�!�;�2�}�W��Y����z��V ��\���u�u�x�<�w�4���������CN�����u�u�u��:�1�4���Y���5��G�����u�u�u�u�w�}�W��Y���@��[�����u�u�&�0�#�/�4���Y����`��C-�����u�u�u�u�w�}�Z����Ʈ�\
��Yd��U���&�=�&��w�}�W���
����V/��N��U���u�u�u�u�z�}��������V�N�����u�|�u�u�w�.����6���F������ �}�g�1� �)�W���B���\��D�����e�1�"�!�w�t�}���:����|��N�����u�|�i�u�8�5����G����]ǑN�U���4�0�!�0���4���Tސ��\��(�����&�8�9�'�6�}����Y����[	��h��3���!�;�=�<�w���������VǻC�����
�u��&�6�)����
����G%��T*������0�3�4�4�4�������OǻC�����
�u��!��1�Ϫ����K��X��ʦ�:�3��u��8����s���E��\1�����4�;�&�4�6�8�8���s���E��\1����� ��u��4�0��ԜY�˺�\	��VN������!�6�u��>����5����F�A�����&�6� ��#�.����6����F��T'����!�u�:�>��<��������A+��F��9�ߊu�u�0�0�>�}����s���F��^��<���4�;�h�u��>�������F�N��Uʷ�:�0�;�u�w�-�������F�N������>�u�u�i�����:���F�N��U���u�u�u�u�w�}�W���Y���F��N�����2�6�u�u�w�.��������F������u�u�u�u�w�}�W���Y���F�N��U���u�u�x�<�w�?�������F��e�����4�6�h�u��<��������JN��X��6����%��9�.�p�F��Y����]F��X���ߊu�u�u��#��W���Y���@"��V#��:���y�u�u�u�w�}�W���Y���F�N��U���u�;�u�<�9�9�F�������9F�N��6���3�;�u�u�j�}�4�������F�N��U���u�u�u�u�w�}�W���Y���K��YN�����1�g�u�:�9�2�W���Yӕ��P��YN��U��u��6�8�9�q�W���Y���F�N��U���u�u�u�u�w�}�ZϷ�Yӕ��]��Y�����:�u�u�u�$�>�������X��v������u�u�u�w�}�W���Y���F�N��U���u�x�:�!�$�:����Nӂ��]��N��Uʦ�6� ��!�4�}�Iϭ�����F��['�U���u�u�u�u�w�}�W���Y���F�N��ʦ�2�0�}�b�3�*��ԶY���p��C�����u��_�u�z�5����Y����G4��V�����6��6�_�w�p����&�Ƨ�Z��~ �����>�4��&�6�>�J�ԜY�˺�\	��VN�����'��9�u��<��������JN��X��6����%��9�.�p�F�ԜY�˺�\	��VN�����4�<�u�'�2�}�Z¨�������R��ʦ�:�3��!�w�p��������w��~ ��1����8� ��w�p��������r��Z'����� ���u�z�+����ӕ��P��B��ʦ�6� ��!�4��W������l��v�����u��6�8�"��Wϓ�����]��NN�����'�6��&�:�1����Y۴��l�N�����6�8�%�}�w�}�Wϵ�����]%��^ ��Kʾ�4��&�4�4�`�^���Tӏ����[�����u�:�!�8�'�u�W���Yӵ��C
��[��U��u�4�%�0�;�q�W���Y���F�N��U���u�u�u�u�w�}�ZϷ�Yӕ��l
��^ךU���u��!��;�9�W��Y����F�N��U���u�u�u�u�w�}�W���Y���F�N�U���u�:�9�4�]�}�W���+����A��[��Kʦ�!�'��9��1�ǵ�����R
��^�����u�u�|�u�z�}��������]l�N�����4�;�u�u�w�c��������F��N��U���u�u�u�u�w�}�W���Y���K�^ �����0�}�b�1� �)�}���Y�ƿ�\��~ ��U���k�&�:�3��)�W���Y���F�N��U���u�u�u�u�w�}�Z����ƿ�T��\����!�_�u�u�w��������[�D/�� ����u�u�u�w�}�W���Y���F�N��U���u�x�u�;�w�4����M�ƨ�D��=N��U����6�8� �w�}�J���8����|��N��U���u�u�u�u�w�}�W���Y���F�C�� ���<�;�1�a�w�2����Y�����T�� ���9�h�u��4�0��������F�N��U���u�u�u�u�w�}�W���TӉ����Y��A���:�;�:�_�w�p�#�������@5��E�����9�,�"�9�w�.���������������:�1�;�u��<��������RǻC����2�'�!�0�4�1��������UF��RN�����4�:�;�u�1�>��������@J��_��U���3�<�<�;�$�}�Z�������V��T�� ���u�;�!�0���W���Y����R��Z�����'�&�9�u�$�/�����Ƹ�Vl�C��4���8� �u� �'�)�������F��T��:���4�<�u�h�$�)��������R��d�����6�0�4�r�>�5�L��Ӵ��l