-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��V�����%�#�1�x�w�(����Y����'��R�����u�'�2�;�;������Ɯ�z��Z������!�o�d�w�(���H���9K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�x�}�~�o�F�������T��y�����u�;�!� �2�)�W���	����Z	��C�����<�=�&��$�/��ԑTӨ��Z	��[N�����8�;�&��#�/��������R��Yd�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Zώ�����	F��V�����<�0�3�'�#�8��������_F��C�����:�{�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���Q��NN��0���"�'�n�u�"�8�>���W����_	��T1�C���9�n�u� �2��2�������P9��S@���ߊu�&�u�:�<���������V��X�����;�&�4�9�]�����Ӷ��u��C'�����<�_�u�x�w�5�W�������R
��Y�����!�'�"�'�$�?�W���������X�����%�9�%�4�2�;����W���F��RN�����4�0�3�9�2�}�ϭ�����JF��Q�����3�'�0�6�w�<����Uӄ��VǻC����=�u�:�'�$�2����Y����V/��:��U���!�'� �0�w�2�W���Ӷ��@��DN�����4�_�u�x�>�)��������	��VN�����<�!�'�&�8�8�W�������JH��XN�����4�0�4�;� �;����s��� �������0�u�=�&��}�ϰ��Ƹ���C�����6�4�4�!�%�.��������G��X�����_�u�x�3�;�8�}���TӲ��$��RN�����u�4�u�0�>�3�ϸ�Ӈ��Z��E�����;�:�u�e�w�3�W�������ǻC����%�4�0�3�;�8�W�������[F��d��X����&��9�2�����?����AF����ʣ�9�1�4�u�g�}����������V�� ���4�2�1�_�w�2����Ӎ��@��[��<���'��6�:�w�}��������W��d��X����9�%�4�2�4����������X ��U���<�u�!�f�w�3�W�������V��YN�����2�1�_�u�8�.��������C��R(�����0�2�=�u�w�3����Y���]ǻ�����!�>�=�&��3����Y����T��S��L�ߊu�:�&�4�#�6��������T��N�����'�o�u�c�]�}�Z����Ư�V ��T��ʶ�9� �4�<�9�)����AӅ��_��9�����u�:�1�9�.�2����
����_ǻC����4�0�#�9�3�9����Ӓ��+����ʺ�u�=�u�4�2�>�����ƫ�GF��RN�����6�0�!�{�w�p�W����Ə�R��Y	��6���3�4�6�<�2�8��������V��_�����!�0�%�%�;�3�W����ƿ�A��B��U���u�:�=�<�w�5�W���5Ӆ��VF��SN��ʙ�7���1�6�/��ԜY����G�������4�6�<�0�2�<�W�������AF��V�U���u�!�!�>�$�)��������@F���� ���:�!�!�0�%�:�Ϻ��ƾ�R��S
�����;�u�0�1�#�8�W��Y����R
��V�����u�=�u�0�8�$�W���Y������D�����4�4�<�u�2�(��������U%��T>�����4�u�u�_�w�p�����ƣ���V�Uʶ�;�!�;�u��)�!�������JF��^ �����o�u��0�1�<��������JF�UךU����u�4�0�w�*�W�������\F��^�����!�0�u�0�3�9��������[��e"�����,�u�:�u�?�.�������K��s��<����<�u�0�6�8�W�������eF��V	��ʷ�u��0�3�6�>��������F��x�����>�6�6�0�y�}�Z���Ӓ����R��ʱ�9�,�'�$�>�8����Y����P��P�����=�u���3�.�������eF��V	�����x�u�:�9�w�8�Ϫ�Y����C��R
�����u�6�;�!�9�}�3���0����V
��T�����0�u�h�>�8�;�4���)����V
��C��N�ߊu�x��!�w�2����Ӓ��5��Q�����!�'�u�;�'�>�����Ƨ�R��R�����9�{��0�;�.�W���s������� ���u�0�0�u�6�<����Y����G	��E��U���u�=�,�4�;�.��������R��T�����:�_�u�x�#�8�ύ�����V��C��[���x�u�4�=�4�<�ϱ�Y����V��Y	�����u�4�u�!�%�}��������R��YN��U���<�3�'�;�]�}�ZϺ��ƿ�^�������&�<�!�'�0�.����s���3��^	��ؔ�'�,�!�u�$�(����Ӗ��C��C�����4�4��1�2�.�8����ƹ�V��YN���ߊu�x�6�9�"�<����������D�����=�u��4�4�0����Ӆ��]��d�����u�;�<�;�3�����ӏ��R��NN�����'�9�'�;�2�c�W�������]��N�����u�|�_�u�z�}��������J����U���4�0�u�0�2�)�W���Ӓ����C��%���'�%�2�!�8�}����T�ƨ�G��Y
�����u�:�0�8�9�:����W����J��g�����<�u�'�4�w�}�����ƾ�]��	N�����;�<�;�1�<�5��������F��@ ��U���_�u�,�0��)�8���ӏ��R��NN�����'�9�'�;�2�c�^ϱ�Y����V��s��:���0�2�=�x�f�9� ���Y����9F�N�����:�3��'�.�>�����ƭ�_F��RN�����9�u�4�0�4�8������������ʘ��u�x�u�2�9�W��� Ӈ��F��CN��U���&�9�&�y�$�3�ϱ�����r%��@��U���0�6�'�u�1�)����T�ƾ�@�u��ʺ�u�=�u��4�3����ӑ��@��T�����<�=�u� �$�)��������P��CךU���3�'�4�%�%�4����Y����R��B��ʡ�0�>�#�'�;�>�1����Ƽ�A��C�����4�u�<� �2�}�Z����Ƹ�VF��P�����;�u�3�6�2�;�����Ʃ�P��E�����2� �<�u�>�1����s�ƪ�]��X �����:�3��4��/�ǵ�����G��RN��U���u�u�;�0�2�f�W���Y���F�N��U���u�u�u�u�w���������P��N��Oʼ�!�2�'�_�w�8����*����r��CU�����4�>�2�u�<���������l��V�����:�,��2�%�>�>����ƥ�9l�Q�����u�4�6�:�1���������~��Y�����u�u�u�u�w�3����B���F�N��U���u�u�u�u�w�}�W���6����_	��q�����u�o�<�!�0�/�}�������5��X�����<�_�u�u�6�4����+����]'��V��U���f��,�!�f�o�W������F��F�����u�k�}�!�2�.�J���I���9F�C�!���u�:�&�4�#�4�W���Y����V��QN�����:�3�<�<�9�.����Y������X������u�0�:�.�4�}���Y����U ��C@ךU���x��#�;�6�>����Ӗ��@�R��U��� �9�6�0�1�>��������_��SN�����0�:�3�0�w�/�ϻ����F������;�u�:�3�>�4���� Ӎ��@��[��<���'��6�:�w�<�Ͻ�����Z��D@��0���u��u� �#�}�W��Y����F
��RN�����9�6��6�8�}��������G��X�����u� �%�!�]�}�W���
������Z,�����3��"��4�}�W�������	[��x�����>�4�!�'�}�6��������z��E�����n�_�u�u�z�	��������]��DN��ʻ�8�0�u�3�5�.�W�������V�������0�u�;�0�4�}�6�������l�N�U���"�u�<�u�8�}�����Ƹ�VF��R��Wʳ�;�!�:�4�>�$�W���Ӈ��[������!�u�u�:�;�}����Y���F��V�����'�;�0�%�6�)�Ϯ�
����VF��D�����<�<�;�&�1�/����Y����R
��X�����;�_�u�u�z�>��������F��Y�����u��u�4�4�1��������P
��\(�����6�0�3�6�2�)�W���Y����	��G�����u�x�!�0�w�6����
����U ��E#��U���9�u�0�0�"�1����6����_	��q�����u��&��;�8�>�������G	��=N��U����!�u�<�4�}�ϭ�	������L�����u� �6�<�9�1�������[����U��� �9�,�&�6�}����Y���F��C��[���=�&�8�4�$�)����ӈ��WF�������;�4�1�!�8�}�5���?����A/��R�����'�7�&�_�w�}�ZϽ�����Z��DN��U���=�8�8�'�y�}�WϽ�����GF��B�����0�3�0��4�}�W�������	[��y�����:�3��"��>�W���;����Z
��E'�����4�!�'�_�w�8��ԜY�ƞ�G��v��¾� ��&��2�;��������\��XN����u�u�u�u�w�}�M���;����\��v�����}�u�>� ��.�4�������~��D��8���;�!�;�0�]�}�W���Y���F�N��U���u�u�u�u�w�}�W�������R��X��%���4�u�u�_�w�}�W���Y���F�N��U���u�u�u�u�w�t�W���Y���F�N��U���u�u�u�u�w�}�W�������9F�N��U���u�u�u�u�w�}�W���Y���F�N��]���8�4�0�:�1�� ������X+��~ �����|�u�u�u�w�}�W���Y���F�N��U���u�|�_�u�w�8����+����]'��V�Uʰ�1��9��2�;��������9��>�����u�:�,��0�/��������9