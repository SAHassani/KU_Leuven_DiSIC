-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B5��q�����=�_�x��#�2�MϚ�Ӥ��VǶN�����4�u�'�?�4�g�'���&����al�*�����c��6�8�2�}�G��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�6�u�g�o�4�������(��^��ʜ�&�'�8�;�$���������9K�v��'���!�u�0�0�!�9�Z�������R
��Y�� ���!�u�;�0�9�1�>�������\ǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x�z�}����
���K�:��ʶ�8�:�0�!�'�)�W���ӣ��R��V��ʡ�2�!�0�u�8�0�����ƣ�G�����߇x�u�>�%�w�(����<����T
��^������u�;�9�3�.��������F
��X��ʡ�0�0�1�:�w�p�W����Ư�R����U���:�;�0�u�1�8�W���Y����^��C�����:�;�u�=�w�/������ƴF�U��[���_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�Զs����R��^��N��� �0�<�0�y�)�(�������R��[�Uʠ�0�<�0�{�"�8�����ȭ�_]Ǒ[�����"�'�n�u�"�8� ���W����BH��[Uװ���!�u�$� ��1����
����V��^��Uʾ�:�3�<�!�w�}�W���Y����]��R��H��n�u�>�4�6�4����Y���	F�������u�h�d�n�w�6��������[F�N����;�0�0�u�j�n�L�������R��R�����o�<�u�;�2�8�W��H��ƹ��TN��U���u�u�u�o�>�}��������W��N�����9�6�u�u�w�}�W�������V��V ��U���:�f�o�u�l�}�������F�N��Oʼ�u�;�0�0�w�`�G���s����l�d�����>�u�u�u�w�}�ϭ�����Z��N������>�-�u�w�}�W���
����\��d�����4�9��!�"��W���ӕ��l
��^�����0��4�w�}�W���Cӏ��@��[���ߊu��0��w�}�W���Y����]F��S1�����_�u��0��3�W���Y�����D�����6�#�6�:�����������Y��E��_�u�&�0�?�4�>���Y�����D�����6�_�u�&�3�/����0���\��YN�����2�6�#�6�8�u�W������]ǑN��1����9�1�;�w�}�W���
����\��d�����!���'�#�}�W���ӵ��w��h��&���d�1�"�!�w�t�}���
����z��T��U���u�;��6�6�<�ǵ�	����W	��C��\�ߊu��!��#�}�W���Y����F��C
�����
�0�!�'�<�(��������F��@ ��U���_�u��!��1����Y���	����*���<�u�n�0�3��$�������lǑV�����!�'�u��w�;�2�������V��DdךU���=�:�
�<�$�<����
����_F��V������!�3�:�m�.��������F��P ��U���4�9��!�"��Mϼ�����l�D�����&�6� ���)�W���&����P9��T��]��1�"�!�u�~�W�W�������@'��B�����u�!�
�:�>�f�Wϭ�����@��T�����o�&�1�9�0�>�}���������D����� �o�&�1�;�:��������Q��X����n�u�&�2�6�}��������F��D�����6�#�6�:��j��������l�C�����&�2�;�_�w�>�����Ƨ�F
��D��U���<�;�1�a�w�2����I������B �����}�g��a�z�����.����O�N�\�ߊu�:�&�4�#�6����
����@��[�����6�:�}�b�3�*����P���V�N�����2�6�#�6�8�u�1���5���F��@ ��U���n�_�u�<�9�1��������G��q����&�1�9�2�4�g�W��B����Z��[N��1����u�u�u�w�}�W���=����GN��G��U���;�:�e�u�j�u����
����G��DS�E���n�_�u�<�9�1��������Z��CN��Oʦ�1�9�2�6�m�}�G��Yӕ��]��D*������9�u�u�w�}��������E��X��:��� ��1�=�f�9� ���Y���F��C����e�|�_�u�>�3�ϭ�����_��B����&�1�9�2�4�g�W��B���T��=N��Xʂ�0�u��6�f�}����Y������D�����&�7�3�9�2�.�Wϛ��ƿ�QK��[��U���&�_�u�x�3�;����ӏ��F�������;�"�<�=�$�?�����ƥ���N�����'�6�&�u�2�8��ԜY����[��X�����;� �&�u�6�8�W�������z��ON��[���"�<�=�&�5�;����Y������d��X���!�4�&�u�2�/��������]��DN��U���!�!�0�3�;�8�ϸ�Ӈ��	��G��U���9�=�#�_�w�p��������Z��Y�����=�u�4�0�8�9��ԜY����[��S��͡� �0�4�,�$�4�ϲ����Y�������u�=�&�;�6�}�����Ƹ�^ǻC�U���u�:�u�-�:�1�W�������J��_��U���9�7�u�:�%�.��������F��RN�����<�9�7�_�w�p��������V��^�����9�u�:�u�6�5�����ƿ�Q ��C��Yʦ�6�u�=�!�>�}��������F������0�9�u�!�#�8������ƹK��N�U���3�9�0�u�w�6����D��ƹK�N��1����}�|�i�w�.��������GN��N��U���x�e�e�8�3�i�J��Y���F��s��<���|�i�u�&�6�<�������F�N��X��d�8�1�a�j�n�W��Y�ƿ�w��~ ��\��u�&�4�4�9�8����K���F�N�Gʸ�1�a�h�g�w�p�W���
����z�N�U���4�4�;�0�8�9�F���Y���F��N����h�d�u�x�w�(����������S��D�ߊu�x�u�&��)�>���P���@��C��3���!�d�u�u�w�}�Z��IӋ��R�_ךU���u�&��!��u�^��Y����G��q����u�u�u�u�z�l�Fϳ����VǻC�Uʦ��!��}�~�a�W�������`��Y
��\���u�u�x�d�e�0���D��ƹK�N��1����}�|�i�w�.��������]�N��U���x�d�f�8�3�i�J��Y���`��^����}��1�-�e�W�W��Yӕ��R��YF�U��&��!���/���Y���F�\��U���u�u�u�_�w�p�Wϭ�=����]N��R�����!���'�#�l�W���Y���T���U���u�_�u�x�w�.�3���0����Z�D������'�!�e�w�}�W���T�����Z��U�ߊu�x�u�&��)�>���P���@��C��&���;�}�|�u�w�}�Z��JӋ��R�]ךU����7�<�!�%�n�_������l�C��U���4�4�;�e�w�`��������Z��]��U���u�x�u�x�w�2�W���Y���K������;�d�u�h�$�����?����T�N��U���u�x�u�:�w�}�W�ԜY�����V����u�h�&��#��1������F�N�U���u�:�u�u�w�W�W��Yӕ��R��YF�U��&��!���/���Y���F�]��U���u�u�u�_�w���������\��N�����&�&��!������Y����G��d�����u�7�2�;�w�}����0ӏ��F������9�:�_�u�w�}�ϗ�D����V��_��U���u�u�&��#��_���E�ƿ�w��~ �����}��1�-��}����*���9F�N�����u�u�u�u�$�����Q���F��s��<���6�;�}�>�9�8�Z�������`��d��U���0�1�<�n�w�}��������9F��Y
�����&�u�;� ��1����B��ƹK��_��*���$�4��4�9�}�2�������]��R �����:�>���4�5����+���F�P�����8�%�}�u�w�}��������[F�N��U���0��1�=�w�}�W��Y���Z��P��O���m�u�u�u�<�<�������F������1�=�u�u�w�p�W���Y����T��S��M���u�u�>� ��>�'��������Z#������2�u�x�w�3�W�������	[�d��U���>�%�u�u�w�}�W���GӍ��PJ�N��U���u�x�u�;�w�3����Y���9F�N��:���6�:�>�u�w�`�W�������P�N��U���<�u�<�!�0�/��������\F��S�����u�:�!�8�'�u�W���Yӵ��C
��[��U���k��8�9��6�W���Y���Z�D�����6�u�u�u��0�������[�d�����>�-�u�u�z�}��������T��N��Uʦ�:�3�:�1�w�}�J���:����\��N��U���u�;�u�!��2��ԜY���@%��Q9��U���u�h�u��2�
�[���Y���K��YN�����:�<�_�u�w�}�4���=���F�
P��6����;�u�u�w�}�ZϷ�Yӕ��l
��^�����'�>�:�3�>�)�Z�������V�N��Uʦ���4�;�9�}�J���
����R��YB��U���u�;�u�!��2��ԜY���@��S�����;�h�u�&�3�/����0���K��YN�����:�<�
�0�#�/�FϺ�����OǻN��U���4�4�4�<��}�Iϭ�=����R
��~ �U���<�u�&�1�;�:����Y����@"��V'��U���u�k�&��#��[���Y���F��N�����4�!�>�%�z�}�������F�N��1���4�'��!�j�}����:����|��N�U���u�!�
�:�>���������W	��C��\��u�u�!�0�$�`�W���Yӕ��P��a�����k�&��6�:�<���Y���\��D�����6�u�u�u�$���������[�D�����9�!�|�u�z�}��������T��S��E�ߠ_�u�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԜY����G����4���8�9�!�'�]�}�Zϊ��ƥ��������6� � �4�8�}����
����F��x�����>�6�6�0�w�2����ӂ��Rl�C�����'�1�6�&�6�.����Y����_�Q�����u�4�%�0�;�}����W�Ƙ�Z��DN�����4�u�x�u��i�W���������^ �����9�8�u�;�w�<�ϭ�����\��NװU���#�:�>�0�����Y����[	��h��3���!�;�=�<�w�<��ԜY�˺�\	��VN����� �4�:�u�%�8�W������l��[�����0�9��_�w�p����&�Ư�N��_��H��r�_�u�x�?�2�(���<����W�N����>�4�6�;�e�z�P���Tސ��\����]���0�&�k�e�~�}�Z¨�������~ ������'�,� �]�}�Z�������P#��I����x�=�:�
�w���������P��N����>�4�6�6�"�}��������FǻC�����
�u���#�2��ԜY�˺�\	��VN�����&�6� ��;�9�W������l��v�����!�u�&�6�"�(����Yӣ��@��OT�����,�"�'�{�&�.�C���+���F�P�����8�%�}�u�w�}����
����[��S����0�u�x�u�9�}�������� ��DךU���u��6�8�;�)����GӒ��VO�C����7�:�0�;�m�}����s���C	����U�ߊu�u�u�9�w�}�W���Y����R��R-��;���u�u�x�<�w�.������ƹF���U���u�u�u�k��)����G���F�N��Uʦ�1�9�2�6�!�>����Nӂ��]��GךU���u���u�w�}�W���^���F�N��U���x�<�u�&�3�1����Y�����v\��U���u�k�r�r�w�}�W���Y���F��N�����2�6�u�u�w�>�W���Y���[������k�e�|�u�z�}��������T��A�����b�1�"�!�w�t�W���YӅ��~F�N��U��r�r�u�u�w�}�W���T�ƥ�F��S1�����u�u�u�6�w�}�W���Y���@��Y�����y�u�x�u�"�}��������E��X��Bʱ�"�!�u�|�w�}�WϽ����F�S����6�8�4�<�{�}�Z����ƿ�W9��P��U���u�6�6�;�w�}�W��Y����C%��E�����x�u�;�u�#�����&����\� N�����u�|�u�u�w�>����Y���[�X��Y���u�u�u�u�z�}��������T��A�����b�1�"�!�w�t�W���YӅ��|��N��U��&��6�8�4�(�[���T�ƣ�GF��S1�����#�6�:�}�n�9� ���Y��ƹF������9�!�u�k�$���������F�N��Uʦ�1�9�2�6�]�}�Zώ�	����"��V8�����!�!�u�4�4�}�W�������	��s=��M�����!�9�m�}��������R��R-��;���u�7�2�;�w�}��������l��RF������>�-�u�?�3�W���Yӕ��R��V��:���i�u�&�6�"�����s���V��^�Uʰ�1�%�:�0�$��8�����ƓF�+��U���������W��Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=dךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Zϑ�-����u ��=N��Xʁ�0�0��r�w�1�ϳ��Ƹ�VF��C�����!�u�=�u�6�-����Y����Z�s(��ʼ�u�u�x�u�$�9��������G��VN�����0�4�9�u�8�}����/Ӡ��rF��D�����=�u�4�4�!�1����T�ƣ�G��N��U���u�&� �0�w�3��������\��B��ʡ�4�&�0�u�%�0�9����״�P
��\d��X���:�4�;�y�6�9��������[��X�����:�u�=�u��.�Wϗ�Y�������� ���;�0�1�u�z�}����Y����_�dךU���4�9��!�"��$���E�Ƣ�GF��^�����!� ��n�]�}�Z�������v��G<�����_�u�x�=�8��W���Y����_��\d��Xǣ�:�>�4�6�4�3����ӕ��P��v�����x�#�:�>�6�>����ӕ��Z��v�����x�#�:�>�6�>����	������V��:��� ���#�w�p��������w��x�����4� ��9�w��3�������A��R �����:�>���'�2����Y۴��l�N�����6�8�%�}�w�}�Wϵ�����QF�N��U���9��7�u�w�}�Z����ƿ�W9��P�����:�}�b�1� �)�W���C�Ɣ�V��^�3�ߊu�u�u��#�(� ������X)��G�����|�u�x�<�w�4������� WǻN�����8�%�}�u�w�}�4���Y���F�	N������>�u�u�w�}�W���Tӏ����h���ߊu�u�u��#��W���Y����@ ��V�����u�u�u�u�z�}��������T��A�����b�1�"�!�w�t�W���YӅ��z��B��U��&��6�8�4�(�[���Y���K��YN�����:�<�
�0�#�/�E�������V�N��Uʶ�;� �%�!�1�`�W�������F��C(�����u�x�<�u�$�9�������F��s��:���u�u�k�&�6�<�������F�N�U���u�!�
�:�>�����ۍ��G��`����1�"�!�u�]�W�W�������F��C(��I����&�7�0�"�-����^����9F�N��ʑ�!��9�1�"�}�ϱ��ƹ�V��X�����!�u�;�0�{�.�W���^�ƻ�@��VN���ߊu�x�3�'�#�8�������t��V�����o�<�u��3�%�GϹ�����VlǻN��X���:�
�u��8��ϑ�����R��V�����u�x�=�:��}�%�������V�N��Xǣ�:�>�4�4�2�8�W���
���F�A�����6�;�&�;�5�8������ƹF������u�9�u�4�'�8��ԜY���E��\1�����&�4�4�4�>�����Y����[	��h��$ʦ�4�4�4�<��)����s���|��B�����9�1�u�;�>�$� ���W����C"��F���ߊu�u�u�0�2�4�W���Y���F�N������9�h�u�g�t�W������G��X	��U��r�r�u�u�w�-�������F�N�����0�u�k�3�;�8�W���Y���F�N�U���u�:�9�4�]�}�W���Y����F�	N�����0� �%�!�1�}�W���Tӏ����[�����u�u�u�9�w�}�J�������p
��N��U���u�u�x�<�w�.������ƹF�N��1���u�h�u�&�6�<����6���F�C����&�1�9�2�4�}�W���YӅ��F�
P��1����9�1� ��1���T�ƣ�GF��S1�����o�u��&�#�<�}�������V��V��2���4�4�4�<�l�W�W�������Z��C"��U��r�r�"�0�w�����D�Ʃ�@��s��#���1� ��9�'�W�Wϭ�����GF�N��U��u��!��#�>�L���
����e��S!��U���i�u��!��1����5����9l��SN��9��