-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s������9�{�=�]�p�6�������\��v�����_�x��<�>�<�W�������6��R1�A߇�x�u�4�0�w�l�=���Y����9K��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�w�>�W��Hӥ��J��_�����;�9��&�%�0����:����A��X חXʔ�9��2�!�w�8�������}��X ��U���!� �0�!�w�3����ӯ��\��C�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z��Y����\��N�����<�0�6�9�"�<�����Ơ�]�������9�!�1�6�2�;�������F�N��U���:�u�4�=���}��T���F�N�����3��8�;�#�3�Ϻ�����]��@��ʶ�0�3�6�0�#�}����
����JF��^חX���u�u�u�u�>�.����W�ƚ�_��A�����4�2�u�'�:�m����W���K�N��U���u�3�&�&��)����Y����@��C��U���;�!�0�4�#�/��������JF����ʳ�'�x�u�u�w�}�W����Ư�V ��T��ʴ�1�1�9�4�;�2�Z���Yӯ��Z��DN�����u�=�;�!�2�0��ԑT���F�N�����<�<�;�u�2�2�Ϸ�Y����l�=C�U���u�u�u��>�}����Ӆ��P��C��ʻ�"�6�0�3�4�8��������P
��\N�����_�x�u�u�w�}�W�������[����ʦ�2�<�<�4�#�-�����ƨ�_��^ �����8�1�9�|�z�W�Z���Y���F��_�����<�<�;�u�6�>����ӏ��R��R��ʷ�u�=�u�:�#�0�F�ԑT���F�N�����0�u�<�&�8�}�'������g��]�����:�3�<�<�9�}�Ϭ��ƣ�Gl�N��U���u�u�3�8�:�/�W�������R��_��Fʷ�!�1�9�4�#�}��������\��^�����x�u�u�u�w�}�W���Y����A��^��ʷ�!�u�3�&�?�.�>����ơ�_��[��U���!�0�d�u�>�W�Z���Y���F��R��U���u�=�;�4�3�9�����ƣ�Z��V�����<�<�;�u�8�>������ƴF�N��U���!�0�9�;�6�}����	����V��X�����;�{�x�_�z�}�W���Y����[��B�����4�1�4�1�"�8�W�������Z��EN�����:�4�<�;�6�8����Y��ƴF�N��U���:�0���o�}��������9K��C��U���u�u�u�=�w�4����ӂ��R��_�����=�&�8�1�;�}�������@HǶd�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�4����Y����F��E�Uʠ�0�<�0�{�#�����&������d�� ���<�0�{� �2�4�(���W����9F��D������2�<�!�;�)����	݇��l�B�����{�>��4�#�2��������\��[�Uʠ�0�"�'�{�<���������U ��^��Ĵ�9�_�x�x�w�$�����Ƹ�R��V������7�4�,��1��������l��U��ʀ���n�u�"�8�"���0�Ț�\��Y��Ĕ��_�x�x�$�3����
Ӓ��]��C�����;�<�,��6�)��������_��Dd�����'�6�_�u�w���������G��RN����2�'�'�;�2�m����P���C	��d��Uʆ�8�9��>�m�4�W���&����P]ǻN�� ���9��0�3�m�4�W�������9F������;�o�<�u�9�4��������R
��_��7���x�u�:�;�8�m�L���Tӳ��W��N�����3��!�o�8�)����������Y��E���u�x�u�g�y�h����?����w��X��6���n�_�'�=�#�>����+����UF��V�����0�3�4�6�>�W�Wϭ�����@+��X��Oʗ��f�
�u�j���������^'��V��6���3�0��&�6�>�^�ԜY����R
��v�����,�o���d��W��>����G%��Q�����'�,�>�:�1���������]ǑN�U���u�=�u�4��)��������F��C�����&�'�u�=�w�4����������[�����=�u�:�3�>�4��ԜY����V��^�����9�6�u��y��W�������GF��G�����u�:�8�0�w�4�����Ƹ�VF��RN�����0�_�u�x�>�}��������^��Z�����;�4�,�:�?�/����Y����V��E�����!�'�7�!�w�<�(�������G��PUךU���'�7�!�u�6�����Y����~��E��U���;�9�<�u�5�2���YӇ��A��C�����!�9�u�3�$�1�:�������@��V�����9�6�w�_�w�.����Y����r
��X��%����o�7�:�2�3�M�������9F��^	��ʦ�&��!�:�1�����Cӄ��_��T�����0�_�u�&�0�<�W�������|��N�����2�6�#�6�8�u�BϺ�����O��N�����u��8�4�6�(�'���Y�ƿ�W9��P�����:�}�`�1� �)�W���s����Z��[N�����8�4�4� �w�}��������E��X��@ʱ�"�!�u�|�]�}����ӕ��G+��s��:���<�0�o�&�3�1��������AN��
�����e�n�_�u�>�3�ϭ�����P��CN����0�}�g�1� �)�W���C����G��DN��U��|�u�x��d�p�}���TӲ����S��Uȸ�u�;�<�0�#�8�3���AӃ��^����U���0�'�&�;�6�4�ϱ�s���5��_�U���6�u�4�u�b�;��������Q��N�����<�<�;�u�2�9�W����ơ�AǻC����!�:�4�u�>�.�����ƥ�G	��_�����0�0�!�!�8�}����ӑ��P��V
�����{�u�6�;�#�3�W�������Z ��N�����9�o�u�n�w�.����Y����U ��[��Oʦ�2�0�}�g�3�*����P���	��R��H���e�|�u�x��n�Z��Yӕ��]��D/��6���3�6�0�!�m�.����Q����\��XN�U��}�!�0�&�j�}�G���Y����U�d�����4�u��!�8�;�3�������Z��SF�U���;�:�e�u�j�u����
���V�N�U��{�d�_�u�$�:����)����z��G�Oʠ�&�2�0�}��0��������Z��]�����:�e�u�h��)����D���O��C��D���_�u�<�;�;�.����0����VW������1�>� ��;�������� F��@ ��U���o�u�:�=�%�}�I���^���F��@�Uʦ�2�4�u��6�8��������F��P ��]���8�4�6�=�$����Jӂ��]��G��H���!�0�&�h�w�m�^���Tӳ��VǑN�����u��0�3�2�)�'���I����Z��SF�U���;�:�e�u�j�u����
���V�N�U��{�d�_�u�$�:����:����Z��Y����o�&�2�0��o��������\������h�u�e�|�w�p�$��T���@��V��6���3�6�0�!�>�8�W�������T��S�����|�o�u�:�?�/�W���^���K�d\�X�ߠu�&�2�4�w����������Y�����3��!�'�9�8�W��Q����A�	N��R��u�x��f�z�W�W�������p	��Q-�����0�o�&�2�2�u�4�������A��RG��H���!�0�&�h�w�m�^���T�Ɵ� H�=d��X���;� �0�!�6�}����,����G%��Q�����&�2�4�&�6�8��������]��^ ��U���u�<�;�9�w�p�W�������[��C�����9�;�u�!�0�.�����ƭ�WF��C�������7�:�<�<�ϰ����F��C�����<�!�u��d�.�WϿ�����G��R��Oʦ�'�;�n�u�6�)����Ӎ��CF��������0�3�<�2�g�����ƥ�D��B�����!�'�7�!�w�8�ϱ�Y����r
��X��%����u�<�;�;�4�Wͪ�����F��C�� ���>�0�u�3�$�5����)����	F��P ��U���w�'�0�n�w�<��������V��X��6���3�0�!��'�m�W�������@F��E��N���4�!�<� �2�6����ӕ��V ��T�����0�o�&�2�6�}�������9F��C�����u�0�%�:�w���������Z��[N��Uȡ� �w�_�u�z�+����
����R��N����>�&�2�;�]�?����s���6��R��ʴ�1�'�%�<�6�8����8����V ��C�����0�3�;�:�#�}��������R��R-��\���7�2�;�u�w�4�W�������W��d�����>�u�=�;�w�}�Wϭ�
����p	��Q>�����h�&�&��#�2���Y�����R/��6���3�<�0�u�j�.��������U]ǻN�����3�_�u�;�w�/����B���K��Y��U���u�:�3�<�>�3�W������ P��UGךU���6�&�}�4�'�8����Yӄ��ZǻN��ʧ�&�;�
�1�2�����:���G��=N��U���x�&�=�&��}�ϻ�����\F��RN������6�8�x�<�2��������]��q������_�u�u�w�p����
����Z��[��ʹ�"�'�!�4�w�m�C�������\��@�����;�0�u�=�w�m�W���Y���_��CN�����<�4�!�<�#�:�ϼ���ƹF������4� �u�h�$�8��������G��EF������}��8�6�>����;���� F��@ ��U���8�4�6�=�$����K���9F�N��8���4�4� ��'�}�Jϭ�����R)��d��Uʰ�1�<�n�u�2�9��������9F�N�����6�0�!�<�w�-����Jӄ��@J��R��U���;�-�u�:�1�4����Y����\��_����_�u��0�1�>����Dӕ��]��D#��1����!�<�0�d�}��������]ǻ�����0�!�u�h�$�:����4����G��C>����u�:�;�:�g�t�}���T�ƅ�U��C�����'�4�0�6�2�;����Ӌ��\��]����u�%�:�0�$�����:���F��P��U���<�u�<�<�0�8��������p
�������u�u�&�9��0���������C#�����!�
�;�0�2�u�'�������}��V������!�x�u�8�3�ϵ�����P6��D�����g�|�n�u�w�}����4����G��C>����u��!�0��)�8���s���V��^�Uʰ�1�%�:�0�$�W�W��Y����U��R �����%�0�u�f�5�)�[Ϛ�����\F��O�����<�<�;�u�$�1� ���H�Ʈ�Gǻ�����3�<�<�;�k�}����ە��G+��s��:���<�0�f�u�8�3���P��ƹ��C-�����9�4�i�u�>�3�ǭ�����w��x�����d�u�:�;�8�m�^�ԶYӖ��P��=�����9�|�u�7�0�3�W����ƾ�@��h���8�9��>�w�5����Y���F��G�����=�u�'�6�>�3�Ϯ��ƣ���V�����0�&�u�=�#�4�W����ƹ���_N��ʶ�'�0�%�;�>�:�W���Y���W��V@ךU���u��4�0�9�4����Dӕ��R��YF�� ���9��4�0�>�.�F�������V�=N��U����4�0�;�>�8�W��
����V/��^��N���u�u�&�=�$��'���K���@6��D��%���d�_�u�u�w�p�4���
�Ʈ�G��YN��ʸ�<�u�:�3�>�4��������R��C�����'�4�0�6�2�;����ӂ��GǻN��U����<�u�<�2�4�ϭ�����F��U�����3�'�!�8�9�}�����Ƹ�VF��v#�����=�u��a��?����Y�����D;��4���:�3��%��}����Y���F��t�����!��%�e�k�}�6�������V
��d��U���0�&�_�u�w�}�W�������_��^��U��&�:�3��;�<�}���Y�Ʃ�WF��d��U���x�u�=�:�2�?����Ӓ����YN�����6�0�!�4�3�)�Ͽ�����G��X�����;�_�u�u�w�p�'�������G��t�����0�!�:�0�2�)�Ͻ�����J�������0�&�!�u�8�}��������^��^�����0�4�_�u�w�}�ǭ�
����p	��Q>�����!�0�_�u�w�}�W�������Z��g��E��u��!�:�1�4����B���F��[��U���u�u�&�:�1�4����)����Z�D-�����<�;�n�u�w�}������ƹF������6�0�!�<�2�}�J���:����Z��Y����_�u�u�;�w�;�}����Ƽ�\��DUװU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�W��s���2��#�����,�1��%�o�}����Y����R��V��U����a��u�8�;����Ӏ����B�����u�x�u�4�3�<�ϸ�����]HǻC�<���&�6�8�4�>�1�W���Ӱ��G��B�����-�c�4�1��/����Y����@HǻC�U���u�;��w�p�W���Y����]F��N�U���u��:�u�]�}�Z���4Ӵ��9F�N��%ʇ�2�u�x�u�w�}�Jϟ�;���F�gN�U���_�u�x�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9F��B�����1��%�m�m�?�������F��Z�����1�%�m�_�w�}�W�������9F�N��U������u�w�}�W���Cӏ��V��T��D�ߊu�u�u�u���3���>���F�T�����0�u�h�d�]�}�W���Y����F�N��U���u�u�u�;�2�8�W��H���F�N��!���������3���:���F�T�����4�u�h����}���Y���r3��e+��!���������(���0�����^ ��O������n�w�}�W���8����f2�N��U���u�o�&�'�9�}�J���0����]ǻN��U�������w�}�W���Y����]��R��H��_�u�u�u�w��0���Y���F�N��U���0�0�u�h�f�W�W���Y�Ǝ�z(��cN��U���u�u�u�u�#�4���YѢ��v%��d��U���u������W���Y���	F��C����u�n�u�u�w�}�4��� ����4��N��U��<�!�2�'�m�}�L���Y���%��pN��U���u�u�u�u�m�4�������]ǻN��U�����u�u�w�}�W���Y����Z��R����u�w�����1���B���F�#��2���u�u�u�u�w�}�MϷ�����\�UךU���u�u� ����>���>���\��Y�����h�d�_�u�w�}�W���6����tF�N��U���u�;�0�0�w�`�F�ԜY���F��c:��;���u�u�u�u�w�}��������\�oL�E��e�e�e�w�]�}�W���Y����F�N��U���u�u�u�;�2�8�W��H���F�N��9����u�u�u�w�}�W�������\�#��>��u�u�u�u���'���<���F�N����;�u�h�w��	�%���s���F�d+��'�����
���}�W������F��r"��4���n�u�u�u�w��:���=���F�N��Oʦ�'�;�u�h�u��2��Y���F��d+�� ���u�u�u�u�w�g��������D��{:��W�ߊu�u�u�u���6���+����g#��T�����2�o�u����3���B���F�;��*����u�u�u�w�}�Mϭ�����	[�x ��M���_�u�u�u�8�)�}���Y���p*��N��U���u�u�u�;�w�)�(�������F�N��4���u�u�u�u�w�}�W���Y����_	��T1�����}�l�1�"�#�}�^�ԜY���F��~ ��U���u�u�u�u�9�}��������E��X��Lʱ�"�!�u�|�]�}�W���Y����gF�N��U���u� �u�!��2��������T��S�����|�_�u�u�w�}�W���Y���F�T�����!�
�:�<��8����H�ƨ�D��^����u�u�u���}�W���Y�������*���<�
�0�!�%�l�W������]ǻN��U���� �u�u�w�}�W������G��X	��*���!�'�d�u�8�3���B���F�-��U���u�u�u�u�m�4�Wϭ�����Z��R����u�:�;�:�g�f�W���Y����F�N��U���u�o�:�!�$�9��������G	��Y�����:�e�n�u�w�}�Wώ�0���F�N��Oʼ�u�&�1�9�0�>����������Y��E��u�u�u�u���#���Y���F��X�����9�2�6�#�4�2�_������\F��d��U���u�����}�W���Y�ƥ�F��S1�����n�u�u�u�w��%���,���F�N��ʦ�1�9�2�6�!�>����Y����G	�UךU���u�u�����>���Y����]F��C
�����6�_�u�u�w�}�6���:����f2�T�� ���!�
�9�2�4�W�W���Y�ƃ�~)��N��U���u�u�;�u�#�����&����\�
�����e�n�u�u�w�}�6���6���F�N����&�1�9�2�4�+����Q�ƨ�D��^����u�u�u����$���Y�������*���<�
�0�!�%�o��������l�N��Uʘ�����w�}�W���ӕ��l��P�����u�u�u� ���9���Y���	����*���2�6�_�u�w�}�W���+����F�N��U���u�!�
�9�0�>�}���Y���f(��e(��"���u�u�u� �w�)�(�������F�N��%��������}�W���Y����F
��^�U���u�u�����2���-����\��D�� ���<�n�u�u�w�}�4���Y���F�N����&�1� �:�>�f�W���Y����v'��N��U���u�o�<�u�$�9������ƹF�N��0�����u�u�w�g����
����_	��TUךU���u�u��d�w�}�W���Y����]F��C
�����6�_�u�u�w�}�2��Y���F�T�����!�
�9�2�4�W�W���Y�Ə�pF�N��U���u�u�;�u�#��������F�N��6�����u�u�w�}��������\��d��U���u����w�}�W���Y�ƥ�F��S1�����n�u�u�u�w��:���Y���F�N��Uʦ�1� �:�<�l�}�W���Yӥ��f*��v<��<���o�<�u�&�3�(����B���F�-��U���u�u�u�u�m�4�Wϭ�����T��=N��U���u���u�w�}�W���Cӏ����h�����_�u�u�u�w��6���8����}F���U���
�9�2�6�]�}�W���Y����3��s+��U���u�;�u�!��1����s���F�e=��U���u�u�u�u�w�3�W���&����Z��N��U�����u�u�w�}�W���Y���@��B����u�u�u�u��	�#���Y���F��^ ����� �:�<�n�w�}�W���+����F�N��U��<�u�&�1�"�2���Y���F��d:��U���u�u�u�o�>�}��������PO��N�����6�8�:�0�#�W�W���
����_F��d��Oʦ�1�9�2�6�!�>����@ӂ��]��G�U���&�2�4�u��1�W�������T��A�����b�1�"�!�w�t�}���Y����R
��t=��U���!�
�:�<��8����M�ƨ�D��^����u�<�;�9�$����
����\��h�����a�u�:�;�8�m�W�ԶYӄ��ZǑN��X���;�!�0���e�[ϟ�������RN��ʥ�%�9�;�u�#�:�W�������[�������<�'�_�u�w�p�#�������GF��#�����;�u�<�0�>�8����ӄ��\��C��%ʴ�1�'�_�u�w�p�#���)Ӕ��F
��^�����!�'�1�7�1�/�W���Y����_F��C��[�ߊu�u�x��$�:�W�������c��N��ʦ�:�3��9�6�4����Ӌ��G��^�����!�{�u�u�$����Y����_	��T1�����}�0�<�0�$�5����)����U��U��Xʆ�e�d�_�u�w�����Dӕ��l
��^�����'�'�&�/����������Z��_�\���x��m�x�]�}�W��Y����T��t�����0�!�<�0�k�j�����ƭ�W��^ ���ߊu�u��9�w�`��������l��C�����/�}��0�1�>����������[�����=�x�>�:�1�����P����V�������=�3�|�u�z��O��s�����V����1�%�m�_�w�}�����ơ�CNǻN��U���&�'�2�h�w�q�W���YӇ��^	��E��H���y�u�u�u�6�8�W���H���F�V�����!�%�!�0�9�9����Y����R
��d��U���4�!�'�&�#�-��������V��X�����k�w���u�W�W���Y����C��
P��1����w�_�u�w�}�������F��=N��U���'�2�h�u�{�}�W�������F�	N��<����y�u�u�w�>��������X�d��U���6�'�,�;�2�/���Y��ƹF�����u�y�u�u�w�0����GӞ�u ��q(��3���y�u�u�u�:�8�W���H���F�Z�����,�;�0�u�i�m�}���Y�ƣ�^	��E��H���y�u�u�u�'�)����D�ƴ�V��^�E��w�_�u�u�w�/���Y��ƹF���*���;�<�2�8�$�}�I���<����`-�=N��U���0�
�4�>�j�}�:���[���F�D�����0�;�h�u��	�2���U���F��D�� ���h�u�����}���Y�ƹ�V9��C�����!�6�u�k�u��'���<����F�N�����8�u�k�w��i�U�ԜY�Ƽ�A��V��U���u�6�>�h�w�<������ƹF���Kʦ��#�_�u�w�}�W���
����l�N����u��9�y�w�}�WϽ�����[�^�����u�u�6�;�j�}�������A��BךU���u�6�;�h�w�2����Y���A�=N��U���6�;�h�u�8�5����G����JǻN��U���'�6�&�<�w�c�P���s���F��[�����u�k�r�r�]�}�W�������X��G�����u�u�6� �w�c����U���F��V�����:�!�h�u�'�3�}���Y�ơ�_��P ����u�%�;�_�w�}�W���Gӕ��_�N��Uʥ�!�0�;�1�#�>�W�������9F�N�����'�1�!�6�w�c����U���F��A�����h�u�%�;�]�}�W�������_	��
P�����_�u�u�u�6�/����D�ƣ�V�N��Uʥ�:�!�h�u�'�3�}���Y�ƣ�^	��S�W��e�e�w�_�w�}�W�������X�^�W�ߊu�u�u�4�%�4����D���V�=N��U���0�d�h�u�f�q�W���YӅ��F�I�Y���u�u�6�4�"�2���Y���9F�N����h�u�d�y�w�}�WϽ����A��d��U���6�6�h�u�f�q�W���YӅ��R��^ ��K��r�_�u�u�w�8�W���^����F�N�����u�k�r�r�]�}�W������A��d��U���6�8�9�6�%�$���Y���9F�N�����h�u�e�y�w�}�WϬ�����\��
P��E���u�u�u�'�#�}�I���^���F�E��U��r�r�_�u�w�}��������J��
P��E���u�u�u�'�#�}�I���^���F�E�����h�u�e�y�w�}�WϬ����A��UװU���x�u�&�<�9�)�Ϛ�)�މ�\��BךU����0�3�4�4�a�W�������c5������� �r�<�=�|�6����*������Y�����3��<�!�~�W�W���Y����XF��[�����1�&�a��]�}�Z�������]��_�� ���!�:�0�8�%�}����YӲ��@F��G�����!�2�u�&�?�/�W�������VF��B�����x�u�0�4�w�8� ���Y����"��V�����>�4�1�!�2��4Ϛ�)�މ�Q
��\d�����0�&��8�;���ԜY����]l�N��U���<�2�0�2��<��������[��N��Uʦ�:�3��9��-�W��
����U%��TUךU���;�u�3�_�w�3�W�������9F�C�����;�:�!� �y�}�W�������GF������4�6�<�0�]�3�W���B�