-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��e�����'�4�{�=�]�p�6�������\��v�����_�x��<�>�<�W�������6��R1�A߇�x�u�4�0�w�e�=���Y����9K��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�w�>�W��Hӥ��J��_�����;�9��&�%�0����:����A��X חXʔ�9��2�!�w�8�������}��X ��U���!� �0�!�w�3����ӯ��\��C�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z��Y����\��N�����'�4�0�u�?�}����Ӌ��G��NN��ʴ�6�8�9�!�w�2�W���Y���F�N��Uʳ�4�!�:�4�w�8�������2����ʼ�&�4�!�4�2�}�W���Mˣ��\��Y��[���x�_�x�u�w�}�W�������G/��_��U��� �1�7�u�%�8��������@F��RN�������<�u�?�}����W��ƴF�N��U����<�u�;�"�8�W���Ӝ��\F��S�����=�u�0� �#�2�W���Y����Z�������u�x�u�u�w�}�W���ӕ��P��YN��6���:�u�=�u��i�2���ӕ��@��C-��ʼ�u�&�0�!�3�}�}��Y���F�:��ʼ�u�0� �'�3�?����Ӿ��Z��[�������3�:�#�3�W�������Z��d�U���u�u�u�u��}�Ϫ�Ӆ��Z�CחX���u�u�u�u�$�>����Ӈ����T�� ���9�4�"�,�w�<�Ϫ�ӕ��VF��[�����x�u�u�u�w�}�W�������GF��Z�����u�=�u�u�"�-�ϱ�Y����w5��+�U���&�&�:�9�w�8�Z���Y���F�B��U���u�=�u�<�6�}����Ӏ��^F��RN��6ʶ�4�;�_�x�z�}�W���Y���@'��B�����u�:�0�u�%�0����)����	��C��1���m�{�u�=�$�.����Y����9K�N��U���u�7�u�:�9�>����ӕ��P��YN��6���:�u�=�u��i�2���Ӓ����CN��6ʼ�u�x�u�u�w�}�W����Ư�R��=C�X���u�u�u�u�w������ƥ�	��NN�����1�<�u��#������ƭ�@��R
�U���_�x�u�u�w�}�WϷ�Yە��@��C-���߇x�u�u�u�w�}�Wϭ�����F�N������u�u�&�6�<����
����U/��=C�U���u�u�u�0�$�W�Z���Y���F������ �u�u��4�0����Yە��G��E��6���3�;�u�u�w�}�}��T���F�N��!���%�%�9�;�w�8��������[F��^�����0�<�u�u�.�1��ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߠ_�<�'�'�w�8��ԜY����Z����*���<�
�d�a�6�1�}���
�ƥ�V��B�����!�{�9�n�w�(�ϩ��Ȝ�T(��C������%�4�9�]�p�Z��� ����@��C�����0�:�3��5�<�φ�����\��^����4�,� ���f����,����~H��X�����&���_�z�p����������Y�����;�_�0�!�#�}����+����C
��z�����_�u�0�0�>�u�W�������G/��_��U���:�9�4�u�l�}����Q���5��G�����u�;�&�1�;�:��ԜY�ƿ�R��V��U���u�;�7�:�2�3�}���Y����G��t��U���;�7�:�0�9�W�W���=����]F�N��U���&�2�0�}�`�9� ���Y����K�d_�D���u�&�:�3��}�W���Y����Z��SF�U���;�:�e�n�w�p�$��HӀ����R��U����f�x�u�8�}��ԜY�ƿ�P��~ ��U���u�;�&�2�2�u�@Ϻ�����O��C�&��l�3�'�<�#�/�[��Y���� F��EN�����u�&�6� ��)�W���Y����@��R
��Bʱ�"�!�u�|�]�}�W�������G*��N��Oʺ�!�&�2�0��j��������]�C��A���u�:�u�;�2�-�W��0��� ��
�����u�'�6��$�0������Ɠ9��_�����0���:�w�/����
����V��TN�����<�;�9�&�2�)�������F������u�h�!� �l�}�����ƿ�]'��B�����u�u�o�7�8�8���Y����l��P�����x��&�1�w�}�$��<Ӆ��U��E�����4���3�9�)��������R��V�����u�=�0�u�9�8����Y���C��[��U���2�&�u� �w�2�W���Y����P	��E��U���6�'�u�7�"�}��������R��S���ߊu�x��<�w�1��������Z��^ ��U���%�3�:�&�8�)��������`6��rN�����0�!�!�u�?�}�������K��^	�����=�!�;�0�w�2����Ӓ����R��ʱ�9�,�:�u�6�<�����ƈ�cHǻ>�����0�0�&�u�5�2�Ϸ�s���@��V��1����9�1�<�2�}�W�������]F�������_�u�u�<�9�1��������W6��R_��U���:�9�4�u�j�)���Y���l�N�����u��&�4�#�<��������Q	��R��O���'�0�_�u�w�p�2����Ƹ�R��_�����<�0�&�2�6�.����Ӓ��G��s=��M���'�u�:�u�2�:�ϩ��ƣ�[��q(��U���x�u�u�0�'�*�Ϯ�Ӊ��@"��V8�����%�e�7�6�"�8��������W6��R_�����2�!�<�2�:�/������ƹF�N�����<�&�4�6�$�2�W���
Ӌ��F
��N�����0�8�1�!�w�8�φ�-ӄ��F��s��#���1�<�0�u�9�W�W���Tӕ��G��[�����u�0�0�7�>�:��������V��DN��U���d�{�u�0�6�.�W���������d��U���u�:�%�9�%�*�ϰ�Ӈ��VF����ʦ�4�4�4�<��-�Fϸ��ƫ�G��PN�����u�<�6�u�#�*����Y���^��^ �����4�4�<��'�m��������UF��RN��9��u��4�u�$�7����Y����A��_�����_�u�u�x��)����Ӎ��CF�������9�1�<�0�w�4�����Ƽ�\��Z@ךU���!�'�7�!�w�8���
����T]ǻN�����7�!�u�0�'�2�W�������Z��G�U���;�9�<�u�#�(�U�ԜY�ƭ�G��B�����u�3�&�4�6�<����	����@��V�����'�0�n�u�w�<��������V��X��'���4�!�4�6�>�8�Mϭ�����Z�C��W�ߠu�7�2�;�w�}�Z��������������0�'�2�&�2�.����Y����\��^
�����=�u��a��}�WϮ�����5��G�����u�u�7�2�9�}�W����ƾ�@��h���8�9��>�w�5����Y�����C�����<�0�u�h�$�<������ƹF�N��1����9�1�<�2�}�Jϭ�����_��^��N���u�u�u�&�2�)��������VV�
N�����'��9�n�w�}�W���Y����F�R �����0�&�_�u�w�p�W�������G��S�����&�2�4�&�4�8�����Ƹ�VF��G�����2�7�:�>�#�}����Y����Z��^��U���&�0�!�'��>����E�ƿ�V��E�����%�e�_�u�w��6�������F�S��1����9�1�<�2�f�Wϻ�ӄ��P��^�����0�&�_�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9F�d��X���=�u�'�6��.��������#��[��U���!�;�<�!�$�<�3���A����\��P��ʳ�'�4���]�}�Zϸ�����]HǻC�<���&�7�!�u�b�<�ψ�Y����R��[�U���u�u�u��8�}�}���T��� ��X �����x�u���0�}�Z���Y�ƞ�Tl�C��U���h���u�z�}�W���Dӫ��UF��R�����6�8�4�1�$�3����+����]��q�����=�<�_�u�z�}�'��Y�͜�z(��QN�����'��6�8�6�9��������V��Y
�����>�<�&���<��ԜY���6�
N��%ʼ�u�;�!�&�2�)�������R��D+������2�u�x�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��N�����0�4�%�0��-�O��������=N��U���%�;�;�u�$�i����Y����V��^��U���u�u�����W���Y���F��^ �����o�u�n�u�w�}�Wϟ�,����a#��N��U���o�<�!�2�%�g�W��Y���F��e+��U���u�u�u�u�w�g�������F��=N��U���u� �����6���+����g#��N��U���o�7�:�0�9�g�W���*��ƹF�N�� �����
����(���<����c2��aN����;�u�h�w���U�ԜY���F��~ ��!���u�u�u�u�w�}�������"��r-��N���u�u�u����2���Y���F�N�����'�o�u�n�w�}�W���;����F�N��U���u�o�<�!�0�/�M���B���F�,��;���u�u�u�u�w�}�Mϭ�����	[�s'��6���_�u�u�u�w��%���+���F�N��U���0�0�u�h�f�W�W���Y�Ə�a4��y=��'���u�u�u�u�9�8����D����F�N��6���u�u�u�u�w�}�W���Y����T��S��N���u�u�u���}�W���Y���F�N�����6�:�u�h��n�1���?����uD��N��U�����u�u�w�}�W���Y����Z��P��O���n�u�u�u�w��;���+����a#��N��Oʼ�!�2�'�o�w�f�W���Y����c+��r<��U���u�u�u�o�>�)����C����9F�N��U�����u�u�w�}�W���Cӄ��l��C��O���w�e�e�e�g�m�G��Y���F��e+��U���u�u�u�u�w�g�������F��=N��U���u��
���}�W���Y�����^ ��O�����w�_�w�}�W���<����g2��yN��U���u�u�!�<�0�g�W͎�-����]ǻN��U����
�����:���Y����G��PN�UȆ����w�]�}�W���Y����~)��N��U���u�u�u�!�>�:�M���*����l�N��Uʀ����u�w�}�W���Y�ƿ�A��T��W�����n�u�w�}�Wϋ�<����g#��h*��0���o�&�'�;�w�`�U���)����gD��N��U��� ����w�}�W���Y����@��Y	��H����a�w�n�w�}�WϮ���ƹF�N��9���u�u�u�u�w�g����
����_	��TUךU���u�u�u�u�w�}�W���Y����]F��C
�����
�0�!�'�e�}�������9F�N��U����u�u�u�w�}�MϷ�Yӕ��l
��^�����'�g�u�:�9�2�G��Y���F��t!��U���u�u�u�o�8�)��������l��C��G���:�;�:�e�l�}�W���YӤ�F�N��U���o�<�u�&�3�1��������AN��
�����e�n�u�u�w�}�5���Y���F�N����&�1�9�2�4�+����Q����\��XN�N���u�u�u���	�W���Y���	F��CN�����2�6�#�6�8�u�@Ϻ�����O��N��U����u�u�u�w�}�W���Y���@��[�����6�:�}�b�3�*����P���F�N��U���u�u�u�u�w�}��������T��A�����b�1�"�!�w�t�}���Y���c%��N��U���u�u�u�;�w�)�(�������P��Z����!�u�|�_�w�}�W���:����F�N��U��� �u�!�
�8�4�(������F��@ ��U���_�u�u�u�w��%���Y���F���U���
�9�2�6�]�}�W���Y����j)��N��U���u� �u�!��2��������U��X����n�u�u�u�w��%���8����F�N��Uʦ�1� �:�<�l�}�W���Yӥ��a?��d-��!���o�:�!�&�3�(����B���F�!��:���u�u�u�u�m�4�Wϭ�����Z��R����1�"�!�u�~�W�W���Y�ƍ�f+��rN��U���u�u�;�u�#�����&����\�
�����e�n�u�u�w�}�4��� ����F�N����&�1�9�2�4�+����Q�ƨ�D��^����u�u�u� ���9���Y�����D�� ���<�n�u�u�w�}�:���*����f2�N����&�1� �:�>�f�W���Y����e#��{!��U���u�o�:�!�$�9������ƹF�N��;�����u�u�w�g����
����_	��TUךU���u�u�����2���-����F��C
�����6�_�u�u�w�}�6���+����v%��T�� ���!�
�9�2�4�W�W���Y�Ə�rW�N��U���u�u�;�u�#��������F�N��4���u�u�u�u�w�}��������\��d��U���u��� ���W���Y�ƥ�F��S1�����n�u�u�u�w��5���Y���F�N��Uʦ�1� �:�<�l�}�W���Yӥ��F�N��U���o�<�u�&�3�(����B���F�-��U���u�u�u�u�m�4�Wϭ�����T��=N��U���u�����}�W���Cӏ����h�����_�u�u�u�w��#���Y���F���U���
�9�2�6�]�}�W���Y����F�N��U���u�;�u�!��1����s���F�t+��9������u�w�3�W���&����Z��N��U�����u�u�w�}�W���Y���@��B����u�u�u�u��	�W���Y���F��^ ����� �:�<�n�w�}�W���+����%��e7��U��<�u�&�1�"�2���Y���F��d:�� ����u�u�o�>�}��������P]ǻN��U�����u�u�w�}�W������G��[���ߊu�u�u�u���W���Y���\��YN�����9�2�6�_�w�}�W���*����F�N��U���;�u�!�
�;�:��ԜY���F��c#��U���u�u�u�u�9�}��������l�N��Uʇ��u�u�u�w�}�W����ƿ�W9��X	��\�ߊu�u�;�u�8�-����B���F��P ��U���-�u�u�!��2��������T��S�����|�_�u�u�>�3�ϭ�	����\��C
�����
�0�!�'�a�9� ���Y����F�D������#�6� �w�.��������V��EF�U���;�:�e�n�w�}�����ƿ�_����*���<�
�0�!�%�i�W������F��NךU���<�_�u�u�z�}�����Ƽ�C��Y�����u�:�!�0��0�����Ƹ�\F��G�����0�4�&�!�w�5�W�����ƹF�N��ʅ�}�0�|�u�2�8������ƹF�N��U���u��a�0�w�}����Y����	�������0�&�4�0�5�;�����Ɓ�^��^�����u�u�x�u�?�}����Ӊ��~F��DN��ʥ�%�9�;�u�#�:�W�������[�������u�u�x�u�?�}�W�������@F��P�����u�0�:�0�#�8����Ӊ��C��=N��U����0�:�8�3�}�����Ɯ�R��EN��ʺ�9�u�0�%�'�1��������_	�������;�!�0�u�w�p�W���M˃�g��R�����!�;�0�&�#�}�Ϯ�	����V��Y�����<�;�9�6�8�6�������K�X�����:�u�=�u��i�Ϫ�Y������B������s��<�'�)����Y����[F��A�����u�x�!�:�4�2�Ͻ�����V
���������m�u�2�2�Ϫ��ƾ�R��C��%ʴ�1�'�_�u�w�p�#�������VF��EN��]����6�8�0�~�>����Y����Z��^ ��U���!�0���o�s�W���Y���g��R��ʡ�0��0�4�;�}����Y����VF��G�����!�:�4�1�#�2��������P��RךU���x�:�!�<�2�2�W���Y������XN�����!� �u�<�?�)�ϟ�_Ӥ��]��
���ߠu�u�&�%�8�8�K���I����W�@��U���&�4�!�6�"�}����?����z��V�����u�x�u�u�w�W�W���Y���F�L�D��d�u�=�;�$�8����8������RN�U���u���~��}�W���Y���F�^�E��w�u�x�u�w�}�W���s�����O��Hʦ�1�9�2�6�!�>����������R����|�n�_�u�w�.�C׻�����@��Rd��Uʲ�;�'�6�8�'�W�W���Y����P��S�D�ߊu�u�u�9�:�9����D����9F�N�����h�u�y�u�w�}��������l��C��*���0�!�h�u�6�.�[���Y����F��R��*���!�'�
�0�2�)�������D��c-��Y���u�u�4�<�'�)�J���=����gD�N��Uʷ�4�6�0�u�i�l�}���Y�Ʈ�V�	N����u�u�
�;�"�}�I���0����JǻN��U���'�<�'�2�j�}�[���Y����R��^ �����u�k�d�_�w�}�W������JǻN��U���>�h�u�w���1���?���9F�N�����h�u�y�u�w�}��������Z��PN��U���u�u�u�:�:�9����D����9F�N�����'�u�k�-�g�m�G��I����l�N�����u�k�d�_�w�}�W���&����W��h����u������}���Y�ƿ�_9��D��K�����y�u�w�}����	����A�	N��4����w�_�u�w�}�������F��b"��&���u�u�u� �2�-��������V��
P��;������y�w�}�Wϫ�����WF�L��0��|�u�u�%�%�}����Y�����S�&���9��>�_�w�}�W���Gӕ��K�N��Uʷ�h�u�!�
�8�4�(�������w��~ �����u�u�u�k��)����D���O�N��Uʶ�'�,�;�h�w�m�[���Y����P��
P�����'�u�k�r�p�q�W���Yӄ��]F�F�����u�k�r�r�{�}�W���	����X��C
�����
�0�!�'�$�>����P���F�T�����6�;�h�u�g�q�W���YӋ��G��Y��H���e�y�u�u�w�<����D�ƣ�V�N��Uʷ�:�!�h�u�'�3�}���Y�Ư�A��V�� ���k�:�0�y�w�}�Wϳ�����]	��S����y�u�u�u�'�`�W�����ƹF������7�0�0�!�j�}����s���F��C�����0�!�h�u�'�3�}���Y�ƣ�V��X��Kʺ�0�y�u�u�w�(�������F��R �U���u�6�'�,�"�}�Iϱ���ƹF��� ���k�&�9��8�)�}���Y�ƣ�^	��S����:�0�_�u�w�}�������D��^�����u�u�4�'�>�.���Y����JǻN��U���d�h�u�d�{�}�W�������X�I�U���u�6�4� �8�8�J���H��ƹF���D��u�d�y�u�w�}����Y���A�N��Uʶ�6�h�u�d�{�}�W�������A��S�R��_�u�u�u�2�}�I���^���F�T�����k�r�r�_�w�}�W���Y����\9��S�������6�8�2�t�}���Y�Ư�^��T�����h�u�d�y�w�}�WϬ����A��d��U���'�!�9�8�3�}�I���^���F�E��U��r�r�_�u�w�}����D���JǻN��U���4�9�4�'�>�}�I���^���F�E��U��r�r�_�u�w�}�������A��d��U���'�!�u�k�p�z�L���Y���F�D/�� ���!�6�u�h�$�:����*����\��d��U���&�6� ��#�a�W�������`
��UךU���u�9�6�u�%�>�%�������w��+������_