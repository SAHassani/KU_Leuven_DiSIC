-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����9�6��%�!�9�Z�������	F��_ �����8�;�4�1��.�W�������K��E������:�0�!�w����MƴƴF��C�D��� �0�g�d�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=C�]���g�d�u�:�.�4��������R
��Y�� ���!�u�:�%�%�)��ԑTӧ��4��_��'���'�0�_�x��)����Y����A��Y��<���'�4�u�;�8�0����s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x��'�8�8�Wϊ��ƪ�_��X�����!�&�!�0�'�2�����Ʈ�\��Q�����3�4�!�:�6�W�Z���Y���F��R�����u� �;�;�w�3�ϸ�
����P
��\N��U���u�0�9�&�:�1�W������F�N��U���:�4�;�u��}����Y����R��X �����4�%�0�9�w�2����Yӯ��K�N��U���u�=�;�8�!�.��������G	��_�����9�u�:�4�9�*�����ơ�_��[�����u�u�u�u�w�+����Ӊ��`��[���߇x�u�u�u�w�}�#���	����@��PN��U���0�<�u�=�w�+����Y����Z��Y
�����!�0�:�!�"�W�Z���Y���F��V�����'�;�3�'�2�}�����Ƹ�VF��Z��6���1�8�<�{�z�W�Z���Y���F��x�����>�4�!�'�>�9����
ӎ����NN�����>�6�6�0�w�5�������F�N��U���:�u�4�=��0�������9K�N��U���u�>�;� ��0��������_��Y
�����=�"�8�;�w�<����Y������^��X���u�u�u�u�w�8����
ӏ��G��D*�����z�u�'�4�$�}�3���0�����������x�u�u�u�w�}�W�������R��YN�����9�u�z�u�6�/�W���Ӄ��^�������4�'�,�<�]�p�W���Y�����D�����u�<�3�'�9�}��������P��R@�����=�&�'�4�8�W�Z���Y���F��~ �����%�0��'�.�1�W����Ƹ���D�����!�4�u�'�2�(�Ϫ�s���F�N��U���0�6�:�>�6�)��ԑT���F�N��Uʁ�<�u�:� �2�.����Y�Ƣ�DF��[�����;�0�0�,�#�0�W�������R��V�����u�u�u�u�w�<����
����GF��[�����6�9� �4�2�)�ϸ�����\��BחX���u�u�u�u�$�>�����ɝ�\��B�����<�u�4�<�w�5�ϭ�����F��[�����'�&�u�� �p�W���Y���F��C��ʦ�<�!�1�<�#�}��������A��D��ʷ�u�&�0�!�9�}�3���0����ZǶN��U���u�u�"�!�w�<��������]F��V�����{�x�_�x�w�}�W���Yӳ����Z>�����6�&�!�u�9�4��������R��E��U����:�0�&�9�}����s���F�N��U���9�7�u�9�4�9�W�������q
��\�����1�!�'�<�2�)�ϭ��ƣ���=C�U���u�u�u�&�#�/�'�������WJ��d�����&�y�&�0�3�9����Y����VF��T�����&�<�2�x�w�}�W���Y�Ʈ�\��@��U���3�'�u�4�4�1����
ӑ��[F��Q�����&�!�<�2�y�	�ϭ��ƣ�9K�N��U���u�&�6� ��)����Y����@'��B�����u�&�4�&�w���������X��^ ��U���=�x�u�u�w�}�W�������@�������4�6�9�!�$�<�W�������V��s��U���%�!�_�x�z�}�W���Y���g��Z�����4�u�0�'�$�<�����ƭ�@��^ �����'�0�0�{�z�}�W���Y���}	����U���1�4�'�8�$�2��������r��Z!��#���1�1�'�;�w�3�W������F�N��U��� �0��&�#�)�W����ƭ�JF��[����� ��!�4�>�s�Z�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����'�'�u�0�2�}����s�ƹ�VF��R�����:�<�
�d�c�<��ԜY����Z�� �����
�!�{�9�l�}��������c��^;�����0��%�4�;�W�W���Y����6��s�����_�u�&�u�8�6�'�������\��s�����'�4�9�_�2�)��������V��X�����:�u�&�u�0�3����s���X(��g��7���>�u�u�;�>�)��������W��XN�O���n�u�u�>�9�(�$�������A%��[��U���<�!�2�'�%�3�������	[�d��Uʾ�#�'�9�6��>����Y�����^ �����'�;�0�g�#�}�W��J��ƹ��CFךU���4�%�0�9�w�}�ϭ�����Z��N��:����>�o�<�w�)�(�����ƹF��b��'���!�o�<�u�8�1���Y����v��C��3���o�<�u�:�;�<�L�ԜY�ƿ�@��C-�����u�;�7�:�2�3�}���Y����@��T�����o�<�u�;�>�3�ǵ�����@��C��U���;�:�e�n�w�p�E���K�����[������;�&�;�w�}�ϫ�
����WN��S�����|�u�x� �y�W�W���
����G6��D�����o�<�u�:�;�<�!����Χ�F��X�����u�u�u�:�9�2�G��Y����`��C>�����u�;��4�2�/�(���7����\��X��U���u�:�;�:�g�f�W���K����9F������1�0�&�o�>�}��������A�������6�9�6�&�f�9� ���Y����K��@����u��!���1����Ǝ�\
��Y8�����>�;� ��:�1����:����K�
�����e�n�u�u�$�<����Y�ƥ�5��Y��M���4�
�}��'�)��������p��RC����!�u�|�u�z��O��Y����w��~ ��Oʼ�u�<�;�1�o�/����Q����F��Z������6�0�d�3�*����P���5��_װU���x�u�9�u�"�-�����ƾ�T��R��U���u�-�:�!�3�)������ƹF��v������9�1�o�8�)�5�������P�������6�9�6�&�f�9� ���Y����F�D/�� ���!�u�u� �w�<����8������Z>�����6�&�d�1� �)�W���Y���`R��d��Uʦ�6� ��!�w�}��������G'��h��;���'�6�9�6�$�l��������]�C��A���_�;�u�'�4���������X2��d�����!�6� �0����������V��X�����:�u�&�u�z�}��������F��EN��U���%�0�u�0�w�$����
Ӂ��R����ʾ�#�'�9�6��>��ԜY����VF��R
�����!�4�u�;�w�<�ϱ�Y����R��R��ʲ�u�;�:�!�2�2����������VN�����u�x�u�=�$�;�����Ư�_��V��U���u� �7�'�8�}��������R��R�����'�1�:�u�?�W�W��6����_��V�����{�u�3�;�#�2�W�������G��N=������%�!�4�'�8�'��� ����	F��C�����0� �;�<�#�:�Ϸ�s�Ʈ�T��N������0�6�:�<�<����G�Ƨ�]��d�����0��6�0�w�5����Y���F��RN�����1�!�u�4�w�8����ӏ��G���� ���4�&�;�9�w������ƨ�G��V�����u�u�0� �9�l�}���Y����9F�N��Xʁ�0�:�9�u�#�8�W���	����WF��D��ʾ�;� ��8�;�.�������R��Y
ךU���u�x�>�#�%�1��������H��YN�����4�0�0�0�w�4�ϭ��Ƹ�^��B��ʢ�_�u�u�u�z�3�����Ƽ�A��R�����0�u�;�!�2�����ӂ��RF��C�U���u�'�!�'�w�f�W�������U]ǻ��U���6�<�;��;��3���8����I��=N��Xʑ�6�4�0�!�2�3����Y����R��[�����9�&�<�u�?�}��������W�����ߊu�:�&�4�#�6��������Z��N�����'�o�u�4�4�>��������VN��Y��&���9�&�0��4�8�L�ԜY����[��R ��ʺ�u�=�u�:�;�*�����ƺ�P��DN��ʶ�'�3�9�,�$�1����W���F��V�����6�=�&�>�!�/����?����AF�N��ʴ�1�:� �%�#�$�϶�
���F��A������6�:�u��s�:���Y����Z
��V�����'�7�1�<�w�5�W�������F���ʠ�0�u�=�&�$�:����s�ƿ�T��������;�u�u�8�1��������X)��E�����6�:�u�:�9�2�G���D�Σ�[��S����0�n�u�&�0�<�W�������J��N�����;�0�!�'�<�+��������G	��N�����u�|�o�u�8�5����GӀ��@�=d�����4�u� �0��.��������\	��V ��Hʡ� �n�_�u�>�3�ϭ�����]��Z��%���u�u�;�<�9�9����)����q��_�����:�e�u�h��)����D���O��C��G���g�u�&�2�6�}�4���:����@+��B�����0�o� �&�0�8�_�������V�S�����'�u�k�r�p�f�W���A��ƹ��Y�����'��4�0�6�4�'���Y�Ǝ�\
��Y8�����>� ��:��2����Y�ƨ�D��^��O���:�=�'�u�i�;����B����Z��[N������4�0�<�2�}�W���
����l��y�����9�6�&�x�f�9� ���Y���F��C����u�:�=�'�w�c�P���P���3��_�Uʦ�2�4�u��#��!�������\��X�����6�:�}��'�)��������p��RN�Dʱ�"�!�u�|�m�}������� ��D����<�;�9�&�6�<��������`��R
�4���,�!�>�;�"�����
����J��_�����:�e�u�h��)����D����G��DN��R��|�u�x��o�l�Wϭ�����@"��V'�����u�u�<�;�3�e����&�Χ�]��d�����0��6�0�f�9� ���Y���F��C����u�:�=�'�w�c�G���B���`W��d�����4�u��4��9�������3��^	��Ӕ�,�!�>� ��2�5�������W	��C��\��u�:�=�'�w�c�_������F�G�U��� �d�d�_�w�4����
����_��R�����o�7�:�0�9�g�W���
��ƓF��P ��U���0��&�!�m�?�������G��d�����4�u� �0��.��������\	��V ��Hʡ� �n�_�u�>�3�ϱ�����]��Z��U���;�<�;�1�<�(�'�������W��X����u�h�}�!�2�.�J���I����K��]�G���&�2�4�u��1�4�������F��RN� ���2�0�}�u�8�3���Y���\��E��K��r�n�u�x�o�e�Wϭ�����\5��E�����4�<�u�u�8�1��������X(��g��7���>�u�u�u�8�3���Y���\��E��Kʳ�9�0�n�u�$�:����*����c��RN�%���0�'�
�}��0��������K�
�����e�u�h�}�#�8���Yۉ��V��
P��E���n�u�x�g�y�o�Wϭ�����\"��V'�����u�u�:�9�6�����Q����F��Z������6�0�x�f�9� ���Y���F��C����u�4�&�|�]�}����Ӊ��G��a�����0�u�:�9�6�����Q����R��E�����u�u�:�;�8�m�L�ԜY����R
��s��<���o��2�0�f�����ۍ��C��V�����'�,�9�x�w�2����I����N��_��U��}�!�0�&�j�z�P���Y����^�=N�����9�:�4�4�9�}�W�������r��N1����� ��8�9�$�8�4�������\��XN�U��}�!�0�&�j�}�������V�U��Xʆ�m�d�u�&�0�<�W�������F��~N�&���0�d��'�.�)��������J5��RN�Dʱ�"�!�u�|�w�p�$��H����Z��[N�����;� �0��m�����H˧��R����1����,�<�0�z�l��������F�=�[�ߊu�<�;�9�8�8��������	F��D�����'�
�}��:�/���������Y��E���h�}�!�0�$�`�WǱ�����X�I��N���u�d�{�d�w�.����Y����r
��X��U���:�9�4�u�j�;����s����Z��[N������!�4�<��-�W�������]0��C������:��:�<�p�W������F��F�����u�k�3�9�2�f�Wϭ�����\'��B�����0�u�u�4�6�(�6���ۍ��^6��T,�����d�1�"�!�w�t�M�������@F�F�����u�k�r�r�~�}�Zύ�L��ƹ��Y����� ��!�<�2�}�W�������A�������6�9�6�&�f�9� ���Y���F��C����u�:�=�'�w�c�P���P���5��^װUʦ�2�4�u��4�0��������_F��D�����6�#�6�:����������X�
�����e�u�h�}�#�8���Y���l�D������6�8� ��1�W�������G'��h��;���'�6�9�6�$�l��������\������h�u�:�=�%�}�I���^����K��[����<�;�9�&�4�(�8������"��V!��4���!�>� ��8�����T�ƨ�D��^��O���:�=�'�u�i�u����
���V�U��Xʆ�`�e�_�u�>�3�ϱ�����z��OT�����;�1�9�2�;�.�Fǵ�����\��V��ñ�"�!�u�|�m�}�������A��UךU���;�9�:�,�4�2�������]��[�����d�>�#�'�;�>�1����Ϩ�D��^����&�2�4�u��>����0�ƈ�G��C/��*����8�'�6�;�>�������\F��d�����4�u��6�:�(�&�������G'��h��;���'�6�9�6�$�l��������l�D������6�8� ��1��������]0��C������:��:�<�p�W������]ǻ�����:�,�6�:�9�����Y����V��=N��X���:�
�<�&�6�)�W������l��R �����x�:�4�4�9�3��������[������� �u�3�f�y���������GF��Y�����u�0�%�u�2�(����T�Ƹ�VF��Z��U���1�&�<�4�>�3�W���Y����\F��\�����;�u�4�<�%�W�W�������VF��O1�����o�&�'�;�l�}����������h�����:�u��!������Cӕ��]��^��C��_�u�!�'�5�)�W���	����G��PUװU���u�=�&�u�>�3�϶��ƭ���GL�����7�!�u�:�2�.��������[��S��ʲ�!�u�x�u�"�6�Ϸ��Ɵ�U��N�����u�0�1�u�8�?�W���ӊ��Z��V�����0�;�!�0�w�p�W���	����XF��SN�����>�1�8�<�$�;�Ϫ�����9F��C�����u�0�%�:�w�����
����@��V�����'�0�n�u�6�)����Ӎ��CF�������;�'�8�;�m�.����Y���G��UךU���'�7�!�u�2�-����:����J��D#�� ���0�u�<�;�;�4�Wͪ�����F��C�� ���>�0�u�3�8�)��������@��V�����'�0�n�u�6�)����Ӎ��CF��������u�<�;�;�4�Wͪ�����F��C�� ���>�0�u�3�8�<����Cӕ��]��^�����w�_�u�!�%�?��������UF��R�����&�o�&�2�6�}�������9F��C�����u�0�%�:�w�����:����	F��P ��U���w�'�0�n�w�<��������V��X��&���!�=�&��;�9�W�������@F��E��N���4�!�<� �2�6����Ӊ��G��a�����<�;�9�<�w�)����s���F��R�����4�u�4�0�6�����Y����Z��RN��U��� �0�!�4�w�5�Ϻ�Ԓ��VǻC����0�u�;�:���E��Y����VF��R
�����0�4�;�u�8�4�W���ӄ��D�������x��0��<�<�ύ�����_��X�����:�u�<�<�0�W�W�������VF��R��ʦ�6� ��!�6�4�;���Y����R
��DN�����n�u�4�!�>�(�ϵ��ƣ���T�� ���9�o�&�2�6�}�������9F��C�����u�0�%�:�w���������b\��^	��ʼ�u�!� �w�]�}�Z���������CN��ʦ�;�u�<�0�>�8�����ƨ���	��U���9�8�;�0�w�4�ύ�5�ƪ�AF��Z�����!�'�7�!�w�8�ϱ�Y����R/��N ��U���;�9�<�u�#�(�U�ԜY����Z��RN�����3�:� �%�#�$��������������_�0�<�_�w�p�;���Ӓ����B�����9�u�;�!�2�����:����\��YN�����u�=�,�4�2�.�������F��RN�����>�1�8�<�y�}�����ƨ�]��XN�����u�=�'�u�$�<��������F���ʷ�!�0�;�!�2�9����
Ӏ����^ �����'�6�&�}�6�-����P����V��=N��U���'�&�;�
�3�8�$�������F��R ךU���u� �0��$�)����E�ƿ�@��R��N���u�u�&�!�%���������Z��S�����'��4�0�6�4�L���Y����w��~ �����<�0�i�u��)�>�������F�N������6�0�0�#�4���Y����@��T�����_�u�u�u��1�4�������F��R>����u��9��4�8�:���
����9F�N��&���!�=�&��'�}�Jϭ�����[��d��U���&�4�4�;�>�8�W��
����z��=N��U����!���'��K���=����]7��N��Uʦ�0�1�1�'�$�����Dӕ��R��S���ߊu�u�u� �2�1�4�������Z�D;��4���:�3�n�u�w�8�Ϸ�B����]��E����_�u�x��#�5����������Y��U���!�0��0��6�������g�������u�:�0�&�%�W�W��������VN��X���<�u�4�=�5�)��������\��YN��ʡ�8�;�{�u�z�}����
����WF��CN��U���%��:�&�6�.�W���
Ӈ��RF��B��U���6�'�;�/�%�)��ԜY����A	��T�����'�&�u�3�#�8����ӏ��G��'��;ʳ�:�u�=�u�$�3��������@��C�����x�:�u�=�w��1���Y����A��E���ߊu�'�6�&��+����P����V��=N��U���'�&�;�
�3�8�8���:���G��=N��U��� �0��&�#�a�W�������V��G�U���u�:�!�'��<�������F��C��%���0�4�<��'�f�W���YӉ��R��Y�����u�h�&�=�$���������C��N��Uʺ�4�6�,�9�$�4�������@%��T-�����<� ��0�>�8�}���Y�ƣ�G��g����u��4�!�?�.�'���B���F��s��<���9�1�i�u��)�>�������C��N��Uʺ�4�4�;�u�j�.��������z]ǻN��U���!���i�w�����)����l�N�����1�1�'�&�w�`��������V��^�����u�u� �0�;�����E�ƿ�@��C-�����%�n�u�u�2�9���YӃ����T��N�ߊu�x��0�#�}����=����]5��TN�����u�=�!�!�;�.����6����_��q�����!�u�4�%�2�}�Z�������A	��C��&���9��>�1�:�4�Y���������������;�u�<�9�1����Y����@l�C�����#�'�9�u�"�-�Ϙ�
ӑ��]F�������=�u�4�4�$�}��������F��CN������>�u�x�w�2����?����V��CN�����!�,�_�u�z�5����Y����P
��\��&���� �!�'�w�p��������|��T�����!�'�>�#�%�1��������F�A�����>�:�;��/�<����[���F�A�����4�0�0�u�6�.�}���T����X9��u��6����8�9��<�}�Z¨�������V����� �%�!��]�}�Z�������\%��Y��&���� �!�u�z�+����Ӊ��F��V��U���;�� �!�6�4�}���T����X9��X,������2��-�w�-����6����_	��^ �����:�;�0�-�w�3��������|��T������;�� �#�/�_���P�����R��U���u�_�u�u�w���������P��S����'�9�6��4�2�[���Tӏ����R	��U��f�u�u�u�<�2��������F�
P��F���u�u�u�u�w�}�W��Y���@��Y	��H���e�_�u�u�8�)����Q���F��e�����u�u�u�u�j�}����U���F�N��X���;�u�:�9�6�W�W���Y����p
��N��U���u�k��8�;�����Y���K�^ �����9�2�6�u�w�}�������F�N��H�����!� ��.�W���Y����]F��X�����h�!� �_�w�}�W�������F�N��U���0��>�w�}�W���Y���Z�D�����6�u�u�u�8�2����Y���F�
P��&���� �!�u�w�}�W������]��Y�����9�&�d�>�!�/����?����AO��=N��U���� �!�4�>�}�W���D�ƣ�J��X��#���1�u�x�u�"�}�������F�X,������2��-�w�c����P���F�N��U���:�!�7�:�2�3�}���TӶ��V
��RN��ʦ�;�u�<�;�;�}�ϳ��Ƹ�^�������!�u�0�!�w�����*����Z��^�����_�u�x�>�!�/����?����AF�N�����y�:� �%�#�$�ϵ�����\��V��ʶ�6�0�{�u�z�}��������\5��T-�����&�;�!�&�9�8�W�������R��R-��U���0�<�8�1�6�8�Ͽ�����]F��p/�����:�1�_�u�z�	��������VF��RN�����:�;��9�3�)�W���Ӈ����N ��ʺ�,�6�:�;�w�2����
����9F��E�����#�'�9�|�w�?����Y����UF��D��*���0��0��<�}����Y���K�d�����>�<�%�!�$�:��������V��C��ʳ�'�!�<�u�?�}��������W	��^ ךU���u�x�4�1�#�8�W�������E��[�����;�u�=�&�:�<�ϑ�������Y��U���9�2�!�u�w�}�Z�������]��A�����;�!�0�&�4�3�W���Ӊ��|��t�����'�4�'�&�9�W�W���Y����W��X�����0�9�u�;�w�8�Ϫ�����R
�������:�>�4�!�%�>����W���F�N��ʸ�9�<�9�u��}��������Z�������0�&�2�4�w�.����*����\�������u�u�u�x�w�3�����ƣ�R��Y=��ʴ�&�'�&�0�8�:�W�������\F��^����� ��8�9�$�8�4������F�N�����=�u�4�4��0���Y���K�c�����u�'�6�&�>�:����Y����R
��X�����u�;�0�"�w�<�ϱ�����e��SN���ߊu�u�u�x�8�<���� ��ƹF�C�!���;� �0�!�2�����:����\��YN�����4�=�#�9�3�2����Y�������� ���4�:�_�u�w�}�Zϩ�Y�����������&�2�4�&�"�4�ϑ�����J��=N��U���x�u�u�u�z�}�����ƭ�W��E�����9� �!�4�2�5� Ϫ�ӵ��PF��P ��ʴ�0�4�&�2�2�}����Y���K�\!�����6��6�:�w�.�D�ԜY���K�N��U���u�u�u�u���(���Y���F�1��*���
�u�u�u�w�}�(���&��ƹF�C�U���%�0�9�u�w�����Y���O9��h1��*���u�u�u�)���(���Y���F��h1��*���_�u�u�u�z�}�W���Y���F�N��U���
�u�u�
�w�}�(���Yӹ��F��hN��U���u�u�
�u�w��W���Y���)��E-��U���u�
�)�u��!�W����ư�l�K1��Uʩ�
�u�)�
�w�!�(���������=N��U���x�u�u�u�w�}�W���Y�Ɠ�l9��h1��*���
�
�
�
���(���&����l9��h1��*���
�
�
�_�w�}�W��Y����P%��a�����_�u�u�u�z�}�W���T����`��t�����u�)�u�u�+�}�WϢ�Y����F����D���u�g�u�u�g�}�W��Y���9F�N��X���u�u�u�u�w�}�W���Y���l9��hN��U���u�u�u�
���W���Y���F��h1�����u�u�x�u��)�>�������W��g-��U���u�
�
�
���(���Y�ư�l9��h1��*���u�u�)�
��W�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��*���u�u�u�u�w�}�W���&���F�C�����4�;�,�6�?�:�^��*����l9��h1��*���
�)�u�u�+��(���&����F���*���u�u�u�x�]�}�W���T���F�N��U���u�u�u�u���(���&���F�1��*���
�
�u�u�w�}�(���&����ll�N��X���:�4�4�;�.�>�G���Y����OF�N��U���)�
�
�)�w�}�W���YӚ��l9��=N��U���x�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w��(���&����F�N��*���
�
�
�_�w�}�W��Y����R/��N �����|�g�����(���&����l9��N��U���u�)�
�
�+�}�W���T���F�C��U���u�u�u�u�w�}�W���Yӹ��l9��h1��U���u�u�
�
���(���Y���l9��h1��*���u�u�u�x�w�2��������V�N��6���u�u�u�u�w�!�(������F�N��*���
�_�u�u�w�p�W���Y���F�N��U���u�u�u�u�w�}�W���Y����l9��h1��*���u�u�u�
���(���s���F�N�����;�,�6�=�0�t�Cύ�:����l9��h1��*���)�u�u�u�w�}����&��ƹF�C�U���u�x�u�u�w�}�W���Y���9��h1��*���
�
�
�_�w�}�W��Y����R/��V��U���u�u�u�u�w�}�W���Y����l9��h1��*���
�
�
�
���(���&����F�N�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�
���(���&����ll�N��X���:�4�4�;�6�4�W���&����l9��h1��*���
�
�
�)�w�}�W���Y���F��h1��*���
�
�u�u�w�p�}���Y���F��V�����<��!�_�w�}�W��Y���F�N��U���u�u�u�u�w�}�W���Y���F��h1�����u�u�x�u�w�}�W���Y�Ɵ�p9��h1��*���
�
�
�
���(���Y�ư�l9��h1��*���
�
�
�
��W�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��*���
�
�
�_�w�}�W��Y���F�N�&���
�
�
�
���(���&����l9��N��U���u�)�
�
���(���&����F�N�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�
���(���s���F�N��U���u�u�a����(���&����l9��h1��*���)�u�u�u�w�}����&����l9��h1��*���u�u�x�_�w�}�W��S���L�D��_�������}�w�]���S���L�D��_�������}�w�]���S���F�N�U���u�u�u�u�w�}�Wρ�&���F�N��U���
�
�u�u�w�}�W���Y����ll�N��X���:� �%�!�.�>�GƁ�Y���O9��h1��*���)�u�u�)���(���&���F��h1��*���
�
�u�u�w�p�W���Y���F�N��U���u�u�u�u�w��(���Y���F�N��*���u�u�u�u�w�}�(���&���F�N��:��� ��;�}�>�5�(���&����l�N��*���
�
�
�
�w�}�W���&����l9��Kd��U���x�u�u�u�w�}�W���Y���F�N��U���
�
�_�u�w�}�Z���8����|��V��U���u�
�
�
��}�W���&����l9��h1��*���
�
�
�
���(���&���F�C��U���u�u�u�u�w�}�W���Y���F�N��U���
�
�
�
���(�ԜY���K�X/�� ���!�4�<��'�}�(���&����l9��KN��U���u�u�u�u�w�!�(���&����l9��h1��U���u�x�u�u�w�}�W���Y���9��h1��*���u�u�u�u���(���Y���F�h1��*���_�u�u�u�z�}��������F��h��U���u�)�
�
���W���Y����l9��h1��	���u�u�u�
���(�ԶY���K�X*�����,�6�8�&�w�)�Ͽ�
����WF��X��U���9�&�!�u�%�)�W���Y����W�������u�u�x�u�?�}��������W	��^ ��ʡ�0��0��<�9����WӲ����U�����,�9�&�'�&�4��ԜY���K��DN�� ���!�u��%�#�<����)����P
��\!�����'��/�{�w�}�Wϱ�����`��R�����4�;�,�6�8�<���� ����Z��N�����u�|�u�u�w�}�W���Y���F�X=�����;��9�1�6�9�_�������]������4�%�0��%�$����6����R'��d��\��u�u�u�:�6�<�������	��Y�� ���_�u�u�u��)�������	��C��&���}��!� ��3�P�������\��XN����u�u�u�u�w�}�W���Y�Σ�J��X��#���1�4�1�:�.�>����Y�Ƨ�E��[��3���:�u�u�|�]�}�W���,����V��g��U��:�&�'�0�2�f�W�������U]ǻ��U���6�&�n�_�w�<��������V��d������!��8�9�8�W�������G��N=����1�"�!�u�w�8�������K�p��U���u�:�!�:�w�4����Y����	��C��&���u�:�"�u�9�*� ���Y����R��Y�����0�_�u�u�z�;�����Ɵ�^��t�����<�{��'�9�}����UӒ����VN�����0�u�0�u�9�)�����Ʈ�9F�C����<�2�/�'�$�}�"���+����	��E������!���9�}�Ͽ�����R��EN�����y�"�<�=�w�}�Z�������@F��RN�����0� �'�1�#�}���������������&�_�u�u�z�����ӂ����V�����4�0�&�!�%�����Y����F��C��%��� �<��;�%�1� ���Y����AǻN��Xʼ�u�:�0�!�6�}����Y����V�V��ʼ�u�&�4�&�%�8�Y���ӑ��_F��Y��U��� �!�9�<�$�}�W��Y����F
��^�����<�<�=�1�~�}�Wϱ�����e��S)���!��8�;�2�t�K�������a��C>��ʺ�u��!���3�_�������J��_��\���;�u��!����������G��N=�����&�4�9�'����������@6��t��ž�6�4�4�'��'�^��Y�ƣ�R��Y'�����~��!��:�3����s���K�t�����4�0�!�0�:�1����Y����V�������4�;�z�u�9�2�ϭ�������V� ���4�u�u�x�w�4�����ƺ�A��YN��U���;�� �!�#�}�����Ƹ�Z��b6�����4�;�;�0�~�W�W���T���F�N��U���u�
�
�
��}�W���Y����l9��h1��U���u�u�u�
���(���Y���5��G�����u�
�)�u�w�}�W���&����l�N��Uʩ�
�
�
�
�w�}�W�������l9��=N��U���u�u�u�u�w�}�W���Y���F��N��*���u�
�u�u��}�Wρ�Y����lF�1��U���
�u�u�x�w��������F��KN��*���u�
�)�u��!�W����ư�l�K1��Uʩ�
�u�)�
�w�!�(���Y���F�N��U���u�u�u�
���(���&����l9��h1��*���
�
�
�
���(���&����l9��=N��U���u��;��#�<�������K��N��X���:�,�6�:�9�}�W���Y���OF�N��U���)�u�u�)�w�}����YӚ�F��N�U���g�u�u�x�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y����l9��h1��*���
�u�u�x�w�2��������WF��h1��*���
�
�
�
���(������F�N��U���u�
�
�
���(���Y���F�C�����4�;�e�u�w�}�Wφ�Y����F��6��	���u�)�u�u�+�}�WϢ�Y����F����-���u�x�u�:�6�<���Y���OF��N��U���)�u�u�)�w�}����YӚ�QF��N��U����u�u��w�}�Z�������z�N��Uʩ�u�u�)�u�w�!�W����Ɣ��TN��Uʶ�u�u�6�u�w��W���!���K������}�|�u�u�+�}�WϢ�Y����F����-���u�1�u�u�3�}�WϺ�Y����F��6ךU���x�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w��(���&����F�N��*���
�
�
�_�w�}�Z���=����]5��TF�����a���
���(���&����OF�N��U���)�
�
�)�w�}�Z�ԜY���F��V�����0�u�u�u�g�}�W��Y���F��\��	���u�)�u�u�+�}�WϢ�Y����F��N��X�ߊu�u�x�u��)�>�������oN��Uʍ�u�u��u�w��W����ư��KN��Uʩ�u�u�)�u�]�}�W��Y����R/��B��]���u��u�u��}�Wφ�Y����F����	���u�)�u�u�+�}�WϢ�Y���F�=N��U����!�u�=�#�)�ϭ��ƣ�	��C��<ń�u�4�u�0�$�<��������G��Z�����:�4�4�;�9�8�[���Y���^����ʡ�0�8�-�;�!�/��������]F��R��ʺ�!�:�u�:�9�.�}���Y����R/��B��<�!��8�;�2�t�W��Y����R/����1����,�<�0�}�.�����Χ�]��d�����0��6�0�<�>��������VO�N����4�;�;�0�~�v�3���4����W��d��Uʺ�4�4�;� �2��3���4����W��N��Hʺ�4�4�;�}������ ����L��Z�����>�;� ��:�1����:������s��4���<�0�u�d�{�2��������KO�*������1�-�n�w�8�Ϲ�����VF��T�����'�0��n�]�}�Zϝ�����G��G�����;�u�9�6�]�}�Z�������u��C*��%����:�>�u�z�+����Ӎ��G��v�����>�6�4�4�%���ԜY�˺�\	��VN�����0�0�u� �2�����Y����[	��h�����0�9�u�#�%�1�}���T����X9��D;��4���:�3�u� �2�1�4��������X��U���4�0�;�'�:�3�W�������P��R ��U���#�:�>�4�$�<��������]��Y��6����6�0��9�.��ԜY�˺�\	��VN������4�0�4�>�}�$�������V0��^
ךU���=�:�
�u��<����
�ƣ�G��g�����x�#�:�>�6�.��������WF��V�����<��!�_�w�p����&�ƿ�R��Y'��1�����-�1�]�}�Z�������@"��V'��U���!���-�3�W�W�������RF��R�����&��u��6�����
�����X��U���6�8� ��;�9��������e��Sd��Xǣ�:�>�4�&�4�(�8���Y����F��C'ךU���=�:�
�u��>����(Ӊ��P��B��Uʓ�4�!�0��8�����CӃ��Z��@��[���6��6�'�4�1����+���F�P�����8�%�}�u�w�}����)����_	��DN��U���8�'�6�9�4�.�W��Y���Z��P��O���_�u�u�u��)�>��� ����[�\!�����'��/�|�w�p��������V��V ��U���:�g�o�u�]�}�W���Ӌ��NǻN��U���0��&�!�w�}�W���Y����f��e�����u�u�u�u�w�p��������RǻN��U���%�0�9�u�w�}�W���Y����E��[�U���u�u�u�u�w�p����
����\��=N��U��� �0�9��2�;�W���Y���	��R/��6���3�u�u�u�w�}�ZϷ�Yӄ��_��=N��U����4�0�;�%�0����Y���	��V�����8�;�y�u�w�}�ZϷ�Yӓ��Z��SF�� ���4�0�<�&�f�9� ���s���F��V�����&�<� ��2�`�W�������_��^ ��:���u�x�u�;�w�3��������\��XN����u�u��4�#�5�������F������=�&��9�3�}�W���Tӏ��$��[��#���:�}��8�%�>����
���F�N������4�0�u�w�}�W��Y����A��V��U���u�u�u�x�w�3�W���
����l��y�����9�6�&�d�3�*�W���Yӕ��R��S�����u�u�u�k�8�8��������F�N��U���<�u� �&�0�8�N���&�Χ�F��X�����x�_�u�u�w�����/����F�N��H����!���;�9����Y���K��YN�����4��6�:������8����I�d��U���&�4�4�;�w�}�W���Y���F��V�����0��u�u�w�}�Z����Ɵ�T��V�����!�>�4�4�9�/�$���T���F��s��<���u�u�u�u�w�}�Iϱ�����~��S?�U���u�u�x�<�w�����H˧��R��������,�<�0�]�}�W���8����|��V��U���u�h�u��4�0�������F�N�U���u�:�9�4��>����7����\��X��X���u�u�u�&�4�(�8���Y���F�S���� ��!�y�w�}�W���Y���\��s��:���'�
�}��:�/�������ǻN��U���6�8� ��w�}�W���Y����r��Z!��$��u�u�u�u�w�p����=����F��N1������:��:�<�p�W�Զs�Ƌ�])��E��1����!�_�u�8�}��������KF�������6�9�6�&�f�9� ���Y�ƫ�]��CךU���x��!�=�#�8��������A	��C��:����>�1�8�>�}�Ϫ��Ƹ�V��E�����#�1�6�'�2�)����Y���Z��_�����0�9�u�:�6�3�}���Y����V��x��6���_�u�u�0�>�W�W���Y����Z��P1�����#�'�9�|�#�8�}���Y���K��D��ʺ�6� ��!�6�4�'���Y����r��Z!��#���1�4�&�'�$�*����Ӓ��9F�N��U���!�'�0�6�8�6����ӑ��W	��C��U���6�0�u�=�w�<�����Ƹ�^��=N��U���u�3�:� �'�)��������F��Y�����|�!�0�_�w�}�W���Y����F��C8�����%�}� ��4�3����E�ƣ�P��x�����}� ��6�9�8�^�ԜY���F��DךU���u�u�u��4�0��������C��B�����0�|�i�u��>����/����c��!��&���;�0�|�:�w���������Z��B�����0�|�_�u�w�}�W���Y����F�N��X���4�6�u�=�w�<�ϱ���������ʺ�6� ��!�6�4�W�������F�N������6�8� ��1�Ǒ�����]��G�����u�u�u�u�w�2����6����C��x�����1�-�u�h�8�>�����΃�G5��~ ����u�u�u�u�w�2����6����C��x�����1�-�u�h�8�>�����΃�G5��~ ����u�u�u�u�2�9���Y����������u�;�u�'�4�.�L�������V��V��2���#�'�9��#���ԶY���p��C�����<�4�u��]�}�Zϊ�����u��E�����!�0�:�!�"�}��������G	��_�����0�9�u�:�6�3����	����]��_�����3�:�u�=�9�4����T�ƥ���"��3���u�<�2�4�w�5�Ϫ�Ӫ��u6�������:�:�&�'�$�)����
����@Hǻ)��&���9��>�4�6�(�M�������F��T'�����;�>� ��8�����T�ƨ�D��^�����4�0�u�u�z�+����Ӣ��\��GN�����<��:�_�w�}�Z�������X4��R����r�u�u�x�!�2��������GF��[��U���x�#�:�>�6�>�ϭ�����F��Dd��U���#�:�>�4��6�$�������9F�C�����
�u��!��)����ۉ��P��B�����<�0��!�'�����P���K��_��*����&�6� ��)����5����F��T'�����u�u��!�6�4�1���CӃ��Z��@��[���:��%�}�#�t�W���YӁ��V����U�ߊu�u�u�u��.����Y���A�C����&�1�9�2�4�g�W��s���F��E�����_�u�u�u�w�����D�ƪ�_��N��U���u�u�u�u�w�}�W���Y���F�N��U���x�u�;�u�8�1��ԜY���F��YN��U��&�;� �%�#��[���Y���F�N��U���u�u�u�u�w�}�W��Y���Q	��R��U���u�u��>�w�}�Iύ�����_�N��U���u�u�u�u�w�}�W���Y���F�N��Xʼ�u�&�1�9�0�>�W���Y����wF�N��U���&�1�:�<����������Z��G�� ���6�;�0�|�{�}�ZϷ�Yӕ��l
��^ךU���u�u��u�w�`�W�������G0��^
���!�%��1�/�t�W���Y���F�N�U���u�!�
�:�>�}�Jϵ���ƹF�N�����u�=�u�<�6�}�1�ԜY�Ƌ�]��C������!��&�]�}�W���Y�ƥ�V��XN������!�6��g�z��������R��N��U���#�:�>�0��1����Y����F��C�����u�u�u�x�!�2��������G0��I����u�u�x�=�8��W���
����R
��=N��U���x�=�:�
�w��W���6����G ��=N��U���x�=�:�
�w�1�W���	����Xl�N��Xǣ�:�>�4�6�w���������V/��B�����0�|�<�_�w�}�W�������RF������� ��9�}�"���������l�N��:��� ��!��8��W�������\��s(�����u�'�9�_�w�}�W�������PF��GN��U���u�u�u�>�2�8�!���D���O�C�����!�
�:�<�w�`�P���Y���F��X�����}�u�u�u�w�}������� ��D�U���u�u�u�u�w�}�W���Y���K�^ �����0�;�u�u�w�}�WϽ����X��r ������&�u�u�w�}�W���Y���F�N��Uʷ�:�0�;�u�w�}�W���:���F�=�����9�y�u�u�w�}�W���Y���F�C����&�1�9�2�4�}�W���Y����wF�N��U���6�8� ��'��8���	����V�^G�U���<�u�&�1�;�:����Y���F��fN��U��u��6�8�"���������z��OG��\��u�x�:�!�$�9�������X4��R���ߊu�u�u�x�?�2�(���?����@��B�����4�9�%�_�w�}�W�������RF��R��#���r�r�u�u�w�p��������a��CN�����u�u�u�x�!�2��������v��C��3���u�u�u�x�!�2����:����R��R-�����u�u�x�=�8��W�������^)��g��$�!�%��1�/�u�^���Y�����X��U���&�6� ��#�>�&Ǒ�����]��F�����u�u� �%�#�<����	����]��NN������:��%��)�^���Y�����R��U���u�_�u�u�w�}�W���
����_F�I�\���x�<�u�&�3�1����C���l�N��Uʥ�'�u�4�u�]�}�W���Y�ƭ�V��S����0�u�u�u�w�}�W���Y���F�N��X���;�u�:�9�6�W�W���Y���P#��N��Kʦ�;� �%�!��q�W���Y���F�N��U���u�;�u�:�;�<�}���Y���F��\N��U���8�9��<�}�W���Y���F�N��U���x�u�;�u�#�����s���F�N��U���u�k�:�6�"������΃�G5��~ �����|�u�x�u�9�}��������F�N��Uʶ�u�u�u�k�$�>��������)��d�����|�<�|�u�z�}��������T��S��'���!�4�_�u�w�3�W�������!��R�����%�!�4�4��f�}���Y����@��YN��ʶ�&�u�=�u�>�<�W����ƣ�G�����ߊu�u��6�:�(�!���۩��`��Y
��\��u�:�7�:�2�3��������e��S"��]����6�;�0�~�f�Wϻ�Ӂ��V��RN�����%�0�9��#���ԶY���r��P �����<�4�u� �'�)�}���8����|��R����� ��!�6��W�W�������G7�
N������!�6��]�3�W���B�