-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��V�����0�3�6�0�#�s��ԑTӧ��[	��$��ʔ�8�'�4�u�9�}����:����]	ǶN�����4�u�'�?�4�g�'���&����al�*�����a��;�u�g�o�Z�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���6�u�e�g��-����Ө��Z	��[N�����8�;�&��%�2�������r
��e�����0�0�#�1�z�}��������]��B�����;�0�;�9��;������ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�x�u�"�-���Y���� ��RN�����;�u�=�u�8�;��������\��@�����4�&�3�9�2�.��������9K�N��U���u�<�u�u�8�-��������*��a'��[�߇x�u�u�u�w�}�#�������U	��C�����,�6�;�4�9�3�W���Y����U��R ��U�����f�
�]�p�W���Y����������;�1�<�u�?�.����WӲ��U��U��U���0�6�u�9�:�3�W�������A��=C�U���u�u�u�=�$�)�Ϯ�����UF��Q�����;�u�=�u�d�0��������Z��CN�����0�'�&�;�]�p�W���Y����������<�;�u�!�2�;�_��W���R��C��D���0�&�&�2�>�4��������R��C��U���u�u�u�u�2�)�WǍ�J����F����U���9�"�;�u�8�;������ƴF�N��U���x�u�u�u�w�}�W�������u��C*��6���3�6�0�!�y�4���������������<�;�&�<�w�5���Y���F�N�����;�u�0�9�4�.����Y����JF����ʶ�1�u�&�;�w�0�W���
Ӈ��RF��^
�����u�u�u�u�w�	�ώ�����VF��E�����:�u�'�!��:����=����V ��T�����<�<�o�x�w�}�W���Y���H�d�����:�%�;�;�$�r��������w��Z��Ń��z�{�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��Ɠ_��V��<���n�u� �0���Y���&����P9��Z����u� �0���s��������WH��[Uװ%���4�0��2�%�>�3�������P��C���ߊu�,�0���n�(���
Ӈ��R�\����!�u�|�:�w�)�(�������P��]����!�u�|�_�w�>�����Ƨ�\��C-�����1�-�:��>��4���Y����T��S��U���x�i��"�$���������\��^��6��u�u�e�u�w�p�K�������p	��Q'�����'�=�&��g�W�W���s�Ư�]��Y��=���0�!�:�3��9����-����r%��N�����'�o�u�u�w�p�K�������p	��Q'�����'�=�&��g�W�W���N���F�A�����&��0�3�9�8�1�������pV�N��N���6�;�!�;�w���������F��u<��F܊�u�h�}�u�w�p�K�������^	��PךU���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��D��d�d�e�d�f�m�F��H����V��_�E��y�_�u�u�f�l�F��I����W��^�D��e�e�d�d�f�m�[�ԜY���W��_�E��d�d�e�d�f�m�G��H����W�d��U���d�d�d�d�f�l�F��H����V��^�D��d�w�u�u�w��F��H����W��_�E��e�e�e�e�f�m�G���Y���D��_�E��d�e�d�e�g�m�F��I����V��L����u�d�d�d�g�l�G��H����W��^�E��d�e�d�y�]�}�W��H����W��^�D��e�d�e�e�g�l�F��I���F�_�D��d�d�e�d�f�m�F��I����W��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�d�d�u�}�W���[����W��^�E��e�e�d�d�g�m�G��I����FǻN��D��d�e�d�d�f�m�F��H����V��^�E��y�_�u�u�f�l�F��H����V��^�D��e�e�e�d�g�l�[�ԜY���W��^�E��d�e�d�e�g�m�G��I����V�d��U���d�d�d�d�g�l�G��I����V��^�D��e�w�u�u�w��F��H����W��_�E��d�e�e�e�f�l�F���Y���D��_�E��e�d�d�d�g�l�F��I����V��L����u�d�d�d�g�l�G��H����V��^�E��e�e�d�y�]�}�W��H����W��^�D��e�e�e�e�g�m�F��H���F�_�D��d�e�e�d�g�l�G��I����V��_�W���u�u�w�d�f�l�F��I����V��^�E��e�e�e�e�u�}�W���[����W��^�E��d�e�e�d�g�m�G��H����FǻN��D��d�e�e�d�f�l�F��H����V��^�D��y�_�u�u�f�l�F��I����W��^�D��e�e�e�e�g�l�[�ԜY���W��^�E��e�e�d�d�g�l�F��H����V�d��U���d�d�d�d�g�m�G��H����W��_�D��d�w�u�u�w��F��H����V��_�E��e�d�d�d�f�m�F���Y���D��_�E��e�e�e�d�f�l�F��H����W��L����u�d�d�d�g�l�G��I����W��_�D��e�e�e�y�]�}�W��H����W��_�E��e�d�d�d�f�l�G��H���F�_�D��d�e�d�e�g�m�G��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�e�d�d�u�}�W���[����W��^�D��d�d�d�e�f�l�F��I����FǻN��D��d�e�d�d�g�m�F��H����W��^�E��y�_�u�u�f�l�F��H����W��_�E��d�d�d�e�f�m�[�ԜY���W��^�E��d�e�d�e�g�l�F��H����W�d��U���d�d�d�d�g�l�F��H����W��_�E��d�w�u�u�w��F��H����W��_�D��d�d�d�d�f�l�F���Y���D��_�E��e�e�d�d�g�l�G��H����W��L����u�d�d�d�g�l�G��H����W��_�D��d�d�d�y�]�}�W��H����W��_�D��d�e�d�d�f�m�F��H���F�_�D��d�d�e�e�f�l�F��H����V��_�W���u�u�w�d�f�l�F��I����W��^�D��d�d�d�e�u�}�W���[����W��_�D��d�d�e�d�f�l�F��H����FǻN��D��d�d�e�e�g�m�G��H����W��_�D��y�_�u�u�f�l�F��I����V��_�E��d�d�e�e�g�l�[�ԜY���W��_�E��d�e�d�e�f�l�F��I����V�d��U���d�d�d�e�g�m�G��H����W��_�E��d�w�u�u�w��F��H����W��_�D��e�d�d�d�g�l�G���Y���D��_�D��e�e�d�e�g�m�G��H����V��L����u�d�d�d�f�m�G��I����W��_�D��d�e�d�y�]�}�W��H����V��_�E��d�d�d�d�f�m�F��I���F�_�D��e�d�e�d�f�m�F��H����V��_�W���u�u�w�d�f�l�G��H����V��_�D��d�e�d�e�u�}�W���[����W��^�D��e�d�e�e�f�l�F��H����FǻN��D��d�d�d�e�f�m�F��I����W��^�E��y�_�u�u�f�l�F��H����V��^�D��d�d�e�e�f�m�[�ԜY���W��_�E��e�e�d�e�f�l�F��I����V�d��U���d�d�d�e�f�m�F��H����W��_�E��d�w�u�u�w��F��H����W��_�E��d�d�d�d�g�m�G���Y���D��_�D��d�e�d�d�g�l�G��H����V��L����u�d�d�d�f�l�F��I����V��_�D��d�d�d�y�]�}�W��H����V��_�E��e�d�d�d�f�l�F��I���F�_�D��d�e�d�e�g�m�F��H����W��_�W���u�u�w�d�f�l�F��I����V��^�D��e�d�d�e�u�}�W���[����W��^�D��d�e�e�e�f�l�G��H����FǻN��D��d�d�e�e�f�l�G��H����W��_�E��y�_�u�u�f�l�F��I����W��^�D��d�d�d�d�g�l�[�ԜY���W��_�D��e�d�e�d�f�l�F��H����W�d��U���d�d�d�d�f�l�F��H����W��_�D��d�w�u�u�w��F��H����V��_�E��d�d�d�e�f�l�F���Y���D��_�D��e�d�e�d�f�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�e�d�y�]�}�W��H����W��_�E��d�e�d�d�f�l�F��I���F�_�D��d�d�e�d�f�l�G��H����W��_�W���u�u�w�d�f�l�F��H����V��^�D��e�d�d�e�u�}�W���[����W��_�D��d�d�e�e�f�l�G��H����FǻN��E��e�e�e�e�g�m�G��I����W��_�D��y�_�u�u�g�m�G��I����W��_�D��d�d�e�e�g�m�[�ԜY���V��^�E��d�d�d�e�f�l�F��I����W�d��U���e�e�e�e�g�m�F��H����W��_�E��d�w�u�u�w��G��I����W��^�D��e�d�d�d�g�m�G���Y���D��^�E��e�d�d�e�f�m�F��H����V��L����u�e�e�e�g�m�G��I����V��_�D��e�e�e�y�]�}�W��I����V��_�E��d�e�d�d�f�m�G��H���F�^�E��e�d�d�e�g�m�F��H����V��^�W���u�u�w�e�g�m�G��I����V��_�D��d�e�d�e�u�}�W���[����V��^�E��e�d�e�d�f�l�F��H����FǻN��E��e�e�d�d�g�m�F��I����W��^�E��y�_�u�u�g�m�G��H����W��_�D��d�d�e�d�f�m�[�ԜY���V��^�E��d�d�e�e�f�l�F��I����V�d��U���e�e�e�e�f�m�F��I����W��_�E��e�w�u�u�w��G��I����W��_�D��d�d�d�d�g�l�F���Y���D��^�E��d�e�e�e�f�m�F��H����W��L����u�e�e�e�g�l�F��I����W��_�D��e�e�d�y�]�}�W��I����W��_�E��d�e�d�d�f�m�G��H���F�^�E��d�e�e�e�g�m�G��H����V��_�W���u�u�w�e�g�m�F��H����V��_�D��d�d�d�e�u�}�W���[����V��^�D��d�e�e�d�f�l�F��H����FǻN��E��e�e�e�d�g�l�F��H����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�e�d�g�m�[�ԜY���V��^�E��e�e�e�e�g�l�F��I����W�d��U���e�e�e�d�f�m�G��I����W��_�D��e�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�G���Y���D��^�E��e�e�e�e�f�l�G��H����W��L����u�e�e�e�g�m�G��H����W��_�D��e�e�e�y�]�}�W��I����V��^�D��d�e�d�d�f�l�G��I���F�^�E��d�d�e�e�g�m�G��H����W��^�W���u�u�w�e�g�m�F��H����W��_�D��d�e�d�e�u�}�W���[����V��_�E��e�d�d�d�f�l�F��I����FǻN��E��e�e�e�d�f�m�G��I����W��^�E��y�_�u�u�g�m�G��H����V��_�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�d�d�e�f�l�F��H����V�d��U���e�e�e�d�g�m�G��I����W��_�E��d�w�u�u�w��G��I����V��^�E��d�d�d�d�f�m�G���Y���D��^�E��e�e�e�e�f�m�F��H����V��L����u�e�e�e�g�l�G��I����W��_�D��e�e�e�y�]�}�W��I����W��^�E��d�d�d�d�f�l�G��I���F�^�E��d�e�d�e�f�m�F��H����W��_�W���u�u�w�e�g�m�F��H����V��_�D��d�d�e�d�u�}�W���[����V��^�D��d�d�d�e�f�l�F��I����FǻN��E��e�e�d�e�f�m�F��H����W��_�E��y�_�u�u�g�m�G��H����V��_�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�d�e�d�g�m�G��I����V�d��U���e�e�e�d�g�l�F��H����V��^�E��d�w�u�u�w��G��I����W��_�D��e�e�e�e�g�m�F���Y���D��^�E��e�d�d�d�f�l�G��I����W��L����u�e�e�e�g�l�G��I����V��^�E��e�d�d�y�]�}�W��I����W��^�E��d�d�e�e�g�m�F��I���F�^�E��d�e�d�d�g�m�G��I����V��_�W���u�u�w�e�g�m�F��H����V��_�E��e�e�e�d�u�}�W���[����V��^�D��e�d�d�d�g�m�G��H����FǻN��E��e�e�d�e�f�l�F��I����V��^�D��y�_�u�u�g�m�G��H����W��_�D��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�d�f�l�F��I����V��^�D��e�w�u�u�w��G��I����W��_�E��d�e�e�e�f�l�G���Y���D��^�E��d�e�d�d�f�l�F��I����W��L����u�e�e�e�g�m�F��H����W��^�E��e�d�d�y�]�}�W��I����V��_�E��d�e�e�e�g�m�F��I���F�^�E��d�d�e�e�f�l�G��I����V��^�W���u�u�w�e�g�m�F��H����V��_�E��e�d�e�e�u�}�W���[����V��_�E��e�e�e�d�g�m�G��I����FǻN��E��e�e�e�e�f�m�G��I����V��_�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�d�g�l�[�ԜY���V��^�E��d�e�e�d�g�m�G��I����W�d��U���e�e�e�d�g�l�F��I����V��^�D��d�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��d�e�e�d�g�l�G��I����V��L����u�e�e�e�g�m�G��I����W��^�E��e�d�d�y�]�}�W��I����V��^�E��e�d�e�e�g�l�G��H���F�^�E��d�e�e�e�f�m�G��I����W��^�W���u�u�w�e�g�m�F��I����W��^�E��e�e�d�d�u�}�W���[����V��_�D��d�e�e�e�g�m�G��H����FǻN��E��e�e�d�d�f�l�G��I����V��^�D��y�_�u�u�g�m�G��H����V��^�E��e�e�d�e�f�m�[�ԜY���V��^�D��e�d�d�d�g�m�G��H����W�d��U���e�e�e�e�f�l�G��I����V��^�E��e�w�u�u�w��G��I����V��_�D��e�e�e�e�g�m�G���Y���D��^�E��d�d�e�e�f�l�F��I����V��L����u�e�e�e�g�l�F��H����W��^�E��d�e�e�y�]�}�W��I����W��_�E��e�d�e�e�g�l�F��H���F�^�E��e�e�d�d�g�m�F��I����W��_�W���u�u�w�e�g�m�G��H����V��_�E��e�e�e�e�u�}�W���[����V��^�D��e�e�e�d�g�m�G��I����FǻN��E��e�e�e�d�f�l�G��H����V��^�D��y�_�u�u�g�m�G��I����W��^�E��e�e�d�d�f�l�[�ԜY���V��^�D��e�d�e�e�g�m�G��H����W�d��U���e�e�e�e�f�l�F��H����V��^�E��e�w�u�u�w��G��I����W��_�E��d�e�e�e�g�m�G���Y���D��^�E��e�d�e�e�f�l�F��I����V��L����u�e�e�e�g�m�F��H����V��^�E��d�d�d�y�]�}�W��I����V��^�D��d�d�e�e�g�l�F��H���F�^�E��e�e�e�e�f�l�F��I����W��_�W���u�u�w�e�g�m�G��H����W��_�E��e�e�e�e�u�}�W���[����V��^�E��d�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�f�l�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�d�d�g�m�[�ԜY���W��_�D��d�d�d�d�g�m�G��H����W�d��U���d�d�d�d�f�m�G��H����V��^�E��e�w�u�u�w��F��H����V��_�D��d�e�e�e�g�l�F���Y���D��_�D��e�d�e�e�g�m�G��I����W��L����u�d�d�d�f�l�G��H����W��^�E��e�d�d�y�]�}�W��H����W��^�E��e�e�e�e�g�l�G��I���F�_�D��d�e�d�e�f�m�G��I����W��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�d�d�u�}�W���[����W��^�D��e�d�d�e�g�m�G��H����FǻN��D��d�d�d�d�g�m�G��I����V��^�D��y�_�u�u�f�l�F��H����W��_�E��e�e�d�e�f�m�[�ԜY���W��_�E��d�d�e�d�f�m�G��H����V�d��U���d�d�d�d�g�m�F��H����V��^�E��d�w�u�u�w��F��H����W��^�D��e�e�e�e�g�m�G���Y���D��_�D��d�e�d�d�g�m�G��I����W��L����u�d�d�d�f�m�F��H����V��^�E��d�d�e�y�]�}�W��H����V��^�D��d�d�e�e�g�m�F��I���F�_�D��d�d�e�e�g�l�F��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�d�d�e�u�}�W���[����W��_�E��d�e�e�d�g�m�G��I����FǻN��D��d�d�e�e�f�l�F��H����V��_�D��y�_�u�u�f�l�F��I����V��_�D��e�e�e�d�g�m�[�ԜY���W��_�E��d�d�e�d�f�m�G��I����V�d��U���d�d�d�d�g�l�G��H����V��^�D��d�w�u�u�w��F��H����W��^�E��e�e�e�e�f�l�G���Y���D��_�D��d�d�d�d�f�l�G��I����W��L����u�d�d�d�f�m�F��I����V��^�E��e�e�e�y�]�}�W��H����V��^�D��d�e�e�e�g�m�G��I���F�_�D��d�e�e�e�g�m�F��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�d�e�d�u�}�W���[����W��^�D��d�e�e�e�g�m�G��I����FǻN��D��d�d�e�e�g�m�F��I����V��^�D��y�_�u�u�f�l�F��I����V��_�D��e�e�e�d�g�l�[�ԜY���W��_�E��d�e�d�e�g�m�G��I����W�d��U���d�d�d�d�g�m�G��H����V��^�E��d�w�u�u�w��F��H����V��^�E��d�e�e�e�g�m�G���Y���D��_�D��e�e�d�d�g�m�F��I����V��L����u�d�d�d�f�m�G��I����W��^�E��d�e�e�y�]�}�W��H����V��^�E��d�e�e�e�g�m�G��I���F�_�D��d�e�e�e�f�m�F��I����V��_�W���u�u�w�d�f�l�F��I����V��_�E��e�e�d�d�u�}�W���[����W��_�D��e�e�e�e�g�m�G��H����FǻN��D��d�d�d�d�f�l�G��I����V��^�D��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�l�[�ԜY���W��_�D��d�d�d�d�g�m�G��I����W�d��U���d�d�d�e�f�l�F��H����W��_�D��d�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�G���Y���D��_�D��d�d�d�d�f�m�F��H����W��L����u�d�d�d�f�l�F��H����V��_�D��d�e�d�y�]�}�W��H����V��^�E��d�d�d�d�f�l�F��H���F�_�D��d�e�e�e�g�l�F��H����W��_�W���u�u�w�d�f�l�F��I����W��^�D��d�d�e�d�u�}�W���[����W��^�E��d�e�e�e�f�l�F��I����FǻN��D��d�d�e�e�g�l�F��H����W��_�D��y�_�u�u�f�l�F��I����W��^�E��d�d�d�e�f�l�[�ԜY���W��_�E��d�e�d�d�g�l�F��H����V�d��U���d�d�d�d�g�m�F��I����W��_�D��d�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�G���Y���D��_�D��e�e�e�d�g�m�F��H����V��L����u�d�d�d�f�m�G��I����W��_�D��e�d�d�y�]�}�W��H����V��_�E��e�e�d�d�f�l�G��H���F�_�D��d�e�e�e�g�m�F��H����W��^�W���u�u�w�d�f�l�F��I����V��^�D��d�d�e�e�u�}�W���[����W��^�D��d�d�d�d�f�l�F��H����FǻN��D��d�d�e�d�f�m�G��H����W��^�D��y�_�u�u�f�l�F��I����V��^�D��d�d�d�d�f�m�[�ԜY���W��_�E��d�e�d�e�g�l�F��H����W�d��U���d�d�d�d�g�l�G��I����W��_�E��e�w�u�u�w��F��H����V��^�E��e�d�d�d�g�l�G���Y���D��_�D��e�e�e�e�f�l�F��H����V��L����u�d�d�d�f�m�G��H����V��_�D��d�d�e�y�]�}�W��H����V��_�D��e�e�d�d�f�l�F��H���F�_�D��d�d�d�d�f�l�F��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��d�e�e�d�u�}�W���[����W��_�E��d�e�e�d�f�l�F��I����FǻN��D��d�d�e�d�g�l�F��I����W��^�E��y�_�u�u�f�l�F��I����V��_�D��d�d�d�d�g�m�[�ԜY���W��_�D��e�e�e�d�g�l�F��H����V�d��U���d�d�d�d�f�l�G��H����W��_�E��d�w�u�u�w��F��H����W��_�E��d�d�d�d�g�l�F���Y���D��_�D��e�e�e�e�g�m�F��H����W��L����u�d�d�d�f�l�G��H����W��_�D��e�d�d�y�]�}�W��H����W��^�D��d�d�d�d�f�l�G��H���F�_�D��d�e�d�e�g�l�G��H����W��_�W���u�u�w�d�f�l�F��H����W��^�D��d�e�d�e�u�}�W���[����W��^�E��e�d�e�e�f�l�F��H����FǻN��D��d�d�d�d�f�l�F��I����W��^�D��y�_�u�u�f�l�F��H����W��_�E��d�d�d�e�f�m�[�ԜY���W��_�E��e�d�e�e�g�l�F��H����V�d��U���d�d�d�d�g�l�F��I����W��_�E��e�w�u�u�w��F��H����V��^�D��e�d�d�d�g�l�G���Y���D��_�D��e�d�e�d�f�l�G��H����W��L����u�d�d�d�f�l�G��H����V��_�D��e�d�e�y�]�}�W��H����W��_�D��d�e�d�d�f�l�G��I���F�_�D��d�d�e�e�g�m�F��H����W��_�W���u�u�w�d�f�l�F��I����V��^�D��d�e�d�e�u�}�W���[����W��_�D��e�e�e�d�f�l�F��H����FǻN��D��d�d�d�d�g�l�G��I����W��^�D��y�_�u�u�f�l�F��H����V��^�E��d�d�d�e�f�m�[�ԜY���V��^�E��e�e�e�e�g�l�F��H����V�d��U���e�e�e�e�g�m�F��I����W��_�E��d�w�u�u�w��G��I����V��^�E��d�d�d�d�g�l�F���Y���D��^�E��e�e�d�e�g�l�F��H����V��L����u�e�e�e�g�m�G��I����V��_�D��d�e�e�y�]�}�W��I����V��_�E��e�d�d�d�f�l�F��H���F�^�E��e�e�e�e�f�l�F��H����W��^�W���u�u�w�e�g�m�G��I����V��^�D��d�e�e�d�u�}�W���[����V��^�D��e�d�d�e�f�l�F��I����FǻN��E��e�e�e�d�g�m�F��H����W��^�D��y�_�u�u�g�m�G��I����W��^�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�d�d�d�f�l�F��H����V�d��U���e�e�e�e�f�m�F��H����W��_�E��d�w�u�u�w��G��I����V��_�D��e�d�d�d�g�l�G���Y���D��^�E��e�d�d�e�g�l�F��H����W��L����u�e�e�e�g�m�G��H����W��_�D��d�e�e�y�]�}�W��I����V��^�D��d�d�d�d�f�l�F��H���F�^�E��e�d�d�d�g�m�F��H����W��_�W���u�u�w�e�g�m�G��I����V��^�D��d�e�d�e�u�}�W���[����V��_�E��d�e�e�d�f�l�F��H����FǻN��E��e�e�e�d�f�m�F��I����W��_�E��y�_�u�u�g�m�G��I����V��_�D��d�d�d�e�g�l�[�ԜY���V��^�D��e�e�d�d�f�l�F��H����V�d��U���e�e�e�e�f�l�F��I����W��_�D��d�w�u�u�w��G��I����W��_�E��e�d�d�d�f�m�G���Y���D��^�E��d�d�d�d�g�l�G��H����V��L����u�e�e�e�g�m�F��I����V��_�D��e�d�d�y�]�}�W��I����W��^�E��d�d�d�d�f�l�G��I���F�^�E��e�e�e�e�f�m�G��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�d�u�}�W���[����V��^�D��d�e�e�d�f�l�F��H����FǻN��E��e�e�d�e�f�l�G��I����W��_�D��y�_�u�u�g�m�G��H����V��_�E��d�d�d�e�f�l�[�ԜY���V��^�E��d�d�e�d�g�l�F��H����V�d��U���e�e�e�e�g�l�G��I����W��_�D��d�w�u�u�w��G��I����W��^�D��e�d�d�d�f�m�F���Y���D��^�E��e�e�e�e�g�l�G��H����V��L����u�e�e�e�g�l�G��I����W��_�D��d�d�e�y�]�}�W��I����W��^�E��d�e�d�d�f�l�F��H���F�^�E��e�e�d�d�f�m�G��H����W��^�W���u�u�w�e�g�m�G��H����W��^�D��d�d�d�d�u�}�W���[����V��^�D��d�d�d�d�f�l�F��H����FǻN��E��e�e�d�e�f�m�G��H����W��_�D��y�_�u�u�g�m�G��H����V��^�D��d�d�d�d�f�l�[�ԜY���V��^�E��e�d�d�d�g�l�F��H����W�d��U���e�e�e�e�g�l�G��H����V��^�E��e�w�u�u�w��G��I����W��_�E��d�e�e�e�g�m�G���Y���D��^�E��e�d�e�d�g�m�G��I����V��L����u�e�e�e�g�l�G��I����V��^�E��e�d�e�y�]�}�W��I����W��_�E��d�d�e�e�g�m�G��H���F�^�E��e�e�d�d�f�m�F��I����V��_�W���u�u�w�e�g�m�G��H����W��^�E��e�e�e�d�u�}�W���[����V��^�E��d�d�d�d�g�m�G��H����FǻN��E��e�e�d�e�g�m�F��H����V��^�E��y�_�u�u�g�m�G��H����W��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��e�d�d�e�f�m�G��I����V�d��U���e�e�e�e�g�l�G��I����V��^�E��e�w�u�u�w��G��I����V��^�D��d�e�e�e�g�l�F���Y���D��^�E��e�d�e�d�g�l�G��I����W��L����u�e�e�e�g�l�G��H����V��^�E��d�e�e�y�]�}�W��I����W��_�E��e�e�e�e�g�m�F��H���F�^�E��e�e�e�d�g�l�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�d�u�}�W���[����V��^�E��d�e�e�d�g�m�G��I����FǻN��E��e�e�e�d�f�l�G��H����V��^�D��y�_�u�u�g�m�G��I����V��_�E��e�e�e�d�f�l�[�ԜY���V��^�D��e�d�e�e�f�m�G��I����V�d��U���e�e�e�e�f�l�F��H����V��^�E��d�w�u�u�w��G��I����W��_�D��d�e�e�e�g�m�F���Y���D��^�E��d�e�e�d�f�l�G��I����W��L����u�e�e�e�g�m�F��I����W��^�E��d�e�d�y�]�}�W��I����V��_�E��e�d�e�e�g�m�F��H���F�^�E��e�d�e�d�f�l�F��I����V��^�W���u�u�w�e�g�m�G��I����V��_�E��e�e�d�d�u�}�W���[����V��_�E��d�e�e�d�g�m�G��H����FǻN��E��e�e�e�e�f�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�d�f�m�[�ԜY���V��^�D��d�e�d�d�g�m�G��I����V�d��U���e�e�e�e�f�l�G��I����V��^�E��e�w�u�u�w��G��I����V��_�E��d�e�e�e�g�l�G���Y���D��^�E��e�d�d�e�f�l�F��I����W��L����u�e�e�e�g�m�G��H����W��^�E��d�d�e�y�]�}�W��I����V��^�D��d�d�e�e�g�m�F��I���F�^�E��e�d�e�e�g�m�F��I����V��_�W���u�u�w�e�g�m�G��H����W��_�E��e�e�d�d�u�}�W���[����V��^�D��d�d�e�e�g�m�G��H����FǻN��E��e�e�e�d�g�m�F��H����V��^�D��y�_�u�u�g�m�G��I����V��_�E��e�e�e�d�f�l�[�ԜY���V��^�E��d�d�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�E��d�w�u�u�w��G��I����V��_�D��e�e�e�e�g�l�F���Y���D��^�E��d�e�e�d�g�l�F��I����W��L����u�e�e�e�g�m�G��I����W��^�E��d�d�d�y�]�}�W��I����V��_�D��d�d�e�e�g�m�F��I���F�^�E��e�e�d�d�g�m�F��I����V��_�W���u�u�w�e�g�m�G��H����W��_�E��e�e�d�d�u�}�W���[����V��^�D��d�d�d�e�g�m�G��H����FǻN��E��e�e�e�e�f�l�F��I����V��^�D��y�_�u�u�g�m�G��I����W��^�D��e�e�e�d�f�m�[�ԜY���V��^�E��e�d�e�d�f�m�G��I����W�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��F��H����W��^�D��d�e�e�e�g�l�G���Y���D��_�D��d�d�e�d�f�m�F��I����W��L����u�d�d�d�f�l�F��I����W��^�E��d�d�e�y�]�}�W��H����W��^�D��d�d�e�e�g�m�F��H���F�_�D��d�d�e�d�g�m�F��I����V��^�W���u�u�w�d�f�l�F��I����W��_�E��e�e�d�d�u�}�W���[����W��_�D��e�e�d�e�g�m�G��H����FǻN��D��d�d�d�d�g�m�F��H����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�d�g�l�[�ԜY���W��_�D��d�e�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�G��I����V��^�E��e�w�u�u�w��F��H����W��^�D��d�e�e�e�g�m�F���Y���D��_�D��e�e�e�d�f�m�F��I����V��L����u�d�d�d�f�l�G��H����V��^�E��d�d�e�y�]�}�W��H����W��^�E��d�e�e�e�g�m�F��I���F�_�D��d�d�e�d�f�l�F��I����V��_�W���u�u�w�d�f�l�F��I����W��_�E��e�e�e�e�u�}�W���[����W��_�D��d�e�d�e�g�m�G��I����FǻN��D��d�d�d�e�g�l�F��I����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�d�g�m�[�ԜY���W��_�D��e�e�e�e�g�m�G��I����W�d��U���d�d�d�d�g�l�F��H����V��^�E��e�w�u�u�w��F��H����W��_�D��d�e�e�e�g�m�G���Y���D��_�D��d�d�e�e�g�l�G��I����W��L����u�d�d�d�f�l�F��H����V��^�E��e�d�d�y�]�}�W��H����W��_�E��d�d�e�e�g�m�G��I���F�_�D��d�e�d�d�g�l�F��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�e�d�e�u�}�W���[����W��^�E��d�e�d�d�g�m�G��H����FǻN��D��d�d�d�d�g�l�F��I����V��^�E��y�_�u�u�f�l�F��H����V��^�D��e�e�e�e�g�m�[�ԜY���W��_�E��e�e�e�d�f�m�G��I����W�d��U���d�d�d�d�g�m�F��I����V��^�E��e�w�u�u�w��F��H����V��^�E��e�e�e�e�g�l�G���Y���D��_�D��d�d�e�e�f�m�F��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�d�e�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��H���F�_�D��d�e�e�e�f�m�G��I����V��_�W���u�u�w�d�f�l�F��I����V��_�E��e�e�e�e�u�}�W���[����W��^�D��e�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��H����V��^�E��y�_�u�u�f�l�F��H����V��^�D��e�e�e�e�g�m�[�ԜY���W��_�E��e�d�e�e�f�m�G��I����W�d��U���d�d�d�d�g�m�G��I����V��^�E��e�w�u�u�w��F��H����V��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�g�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�e�y�]�}�W��H����W��_�E��d�d�d�d�f�l�F��H���F�_�D��d�e�e�e�g�l�G��H����W��_�W���u�u�w�d�f�l�F��I����W��^�D��d�d�d�e�u�}�W���[����W��^�D��d�e�e�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��H����W��_�E��y�_�u�u�f�l�F��H����V��_�E��d�d�d�d�g�m�[�ԜY���W��_�E��d�d�d�d�f�l�F��H����V�d��U���d�d�d�d�g�m�F��H����W��_�D��e�w�u�u�w��F��H����V��_�E��d�d�d�d�f�l�G���Y���D��_�D��d�e�e�d�g�m�F��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�d�y�]�}�W��H����W��^�D��d�e�d�d�f�l�F��H���F�_�D��d�e�d�d�g�l�G��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��d�d�e�d�u�}�W���[����W��^�E��d�d�e�d�f�l�F��I����FǻN��D��d�d�d�d�f�m�G��H����W��_�D��y�_�u�u�f�l�F��H����V��^�E��d�d�d�d�f�m�[�ԜY���W��_�E��e�d�d�e�g�l�F��H����V�d��U���d�d�d�d�g�l�F��H����W��_�D��e�w�u�u�w��F��H����W��^�D��d�d�d�d�f�m�F���Y���D��_�D��e�e�e�e�g�m�F��H����V��L����u�d�d�d�f�l�G��I����W��_�D��d�e�e�y�]�}�W��H����W��^�D��e�e�d�d�f�l�F��I���F�_�D��d�d�e�d�f�l�F��H����W��^�W���u�u�w�d�f�l�F��I����V��_�D��d�d�e�e�u�}�W���[����W��_�D��e�e�e�e�f�l�F��I����FǻN��D��d�d�d�e�f�l�F��I����W��_�E��y�_�u�u�f�l�F��H����V��^�E��d�d�d�d�g�l�[�ԜY���W��_�D��d�e�d�e�g�l�F��H����V�d��U���d�d�d�d�f�l�G��I����W��_�D��e�w�u�u�w��F��H����W��^�D��e�d�d�d�f�m�G���Y���D��_�D��e�e�e�d�g�m�F��H����V��L����u�d�d�d�f�l�G��H����W��_�D��d�e�e�y�]�}�W��H����W��_�E��d�e�d�d�f�l�F��I���F�_�D��d�d�d�e�g�l�G��H����W��_�W���u�u�w�d�f�l�F��H����V��^�D��d�d�d�d�u�}�W���[����W��_�D��e�e�d�e�f�l�F��H����FǻN��D��d�d�d�d�g�m�G��I����W��_�D��y�_�u�u�f�l�F��H����W��^�E��d�d�d�e�f�l�[�ԜY���W��_�D��d�d�d�e�f�l�F��H����W�d��U���d�d�d�d�f�m�F��I����W��_�D��d�w�u�u�w��F��H����V��_�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�d�d�f�m�G��H����W��L����u�d�d�d�f�l�F��I����W��_�D��e�d�d�y�]�}�W��H����W��_�D��e�e�d�d�f�l�G��H���F�_�D��d�d�d�e�f�l�F��H����W��_�W���u�u�w�d�f�l�F��H����V��^�D��d�d�e�e�u�}�W���[����W��_�E��e�e�d�d�f�l�F��I����FǻN��D��d�d�d�d�f�m�G��I����W��_�E��y�_�u�u�f�l�F��H����W��^�E��d�d�d�d�g�m�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��I����W��_�D��e�w�u�u�w��G��I����V��^�E��e�d�d�d�f�m�G���Y���D��^�E��e�e�e�d�f�l�G��H����V��L����u�e�e�e�g�m�G��H����V��_�D��d�e�d�y�]�}�W��I����V��^�D��e�d�d�d�f�l�F��H���F�^�E��e�e�e�d�f�m�G��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�e�d�u�}�W���[����V��^�D��e�e�e�d�f�l�F��I����FǻN��E��e�e�e�e�f�m�F��H����W��_�E��y�_�u�u�g�m�G��I����W��^�E��d�d�d�d�g�m�[�ԜY���V��^�E��e�e�e�e�g�l�F��H����W�d��U���e�e�e�e�g�l�G��H����W��_�D��d�w�u�u�w��G��I����W��_�E��d�d�d�d�f�m�F���Y���D��^�E��e�e�e�d�f�m�G��H����V��L����u�e�e�e�g�m�G��H����V��_�D��d�d�e�y�]�}�W��I����V��^�D��d�d�d�d�f�l�F��I���F�^�E��e�e�d�e�f�l�G��H����W��_�W���u�u�w�e�g�m�G��H����V��_�D��d�d�e�e�u�}�W���[����V��^�D��d�d�d�e�f�l�F��I����FǻN��E��e�e�e�e�f�m�G��I����W��_�D��y�_�u�u�g�m�G��I����W��_�E��d�d�d�d�f�m�[�ԜY���V��^�E��d�d�e�d�g�l�F��H����W�d��U���e�e�e�e�g�m�G��I����W��_�D��d�w�u�u�w��G��I����V��_�E��e�d�d�d�f�m�F���Y���D��^�E��d�e�d�d�g�m�F��H����W��L����u�e�e�e�g�m�F��H����W��_�D��d�e�e�y�]�}�W��I����V��^�E��d�e�d�d�f�l�F��H���F�^�E��e�e�e�d�f�m�F��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�e�u�}�W���[����V��^�E��e�d�e�d�f�l�F��H����FǻN��E��e�e�e�d�g�l�F��H����W��_�E��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�g�l�[�ԜY���V��^�E��e�d�e�d�f�l�F��H����W�d��U���e�e�e�e�g�m�G��H����W��_�D��d�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�G���Y���D��^�E��d�d�d�d�g�m�F��H����W��L����u�e�e�e�g�m�F��H����W��_�D��d�d�d�y�]�}�W��I����V��_�D��e�e�d�d�f�l�F��H���F�^�E��e�e�e�e�f�l�F��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�d�d�d�u�}�W���[����V��^�D��e�e�e�e�f�l�F��H����FǻN��E��e�e�e�d�f�m�G��H����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�e�e�e�f�l�F��H����W�d��U���e�e�e�e�g�m�F��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�G���Y���D��^�E��d�d�e�d�g�l�F��I����V��L����u�e�e�e�g�m�F��I����W��^�E��e�e�d�y�]�}�W��I����V��_�E��d�e�e�e�g�m�G��H���F�^�E��e�e�e�d�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����W��_�E��e�e�e�d�u�}�W���[����V��^�D��d�e�e�e�g�m�G��I����FǻN��E��e�e�e�d�f�l�G��H����V��^�E��y�_�u�u�g�m�G��I����W��^�D��e�e�e�e�g�l�[�ԜY���V��^�E��e�e�d�d�f�m�G��I����W�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��_�E��d�e�e�e�g�m�G���Y���D��^�E��d�d�e�d�f�l�F��I����V��L����u�e�e�e�g�m�F��I����V��^�E��e�d�e�y�]�}�W��I����V��^�D��d�e�e�e�g�m�G��H���F�^�E��e�e�e�d�f�m�F��I����V��_�W���u�u�w�e�g�m�G��I����V��_�E��e�e�e�e�u�}�W���[����V��^�E��d�e�d�d�g�m�G��I����FǻN��E��e�e�e�d�g�m�G��I����V��^�D��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�f�m�[�ԜY���V��^�E��e�d�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��H����V��^�E��d�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�F���Y���D��^�E��d�e�e�e�f�l�G��I����V��L����u�e�e�e�g�m�F��I����W��^�E��e�d�d�y�]�}�W��I����V��_�D��e�d�e�e�g�m�G��H���F�^�E��e�e�d�d�g�l�F��I����V��_�W���u�u�w�e�g�m�G��H����V��_�E��e�e�e�d�u�}�W���[����V��^�D��d�e�d�d�g�m�G��H����FǻN��E��e�e�e�e�f�l�F��I����V��^�E��y�_�u�u�g�m�G��I����W��_�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�d�e�e�f�m�G��I����V�d��U���e�e�e�e�g�l�G��I����V��^�E��e�w�u�u�w��G��I����W��_�D��e�e�e�e�g�l�G���Y���D��^�E��e�e�d�d�f�m�G��I����W��L����u�e�e�e�g�m�G��I����W��^�E��e�e�e�y�]�}�W��I����V��^�E��e�d�e�e�g�m�G��I���F�^�E��e�e�d�e�f�m�G��I����V��^�W���u�u�w�e�g�m�G��H����W��_�E��e�e�d�e�u�}�W���[����V��^�E��e�d�d�e�g�m�G��H����FǻN��E��e�e�e�e�g�m�G��H����V��^�E��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��d�e�e�d�f�m�G��I����V�d��U���e�e�e�e�g�m�F��I����V��^�E��e�w�u�u�w��G��I����V��^�E��d�e�e�e�g�l�G���Y���D��^�E��e�d�d�e�g�m�G��I����W��L����u�e�e�e�g�m�G��H����V��^�E��e�e�e�y�]�}�W��I����V��_�E��d�e�e�e�g�m�G��I���F�^�E��e�e�e�d�f�l�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�e�u�}�W���[����V��^�E��d�d�e�e�g�m�G��H����FǻN��E��e�e�e�e�g�m�F��I����V��^�E��y�_�u�u�g�m�G��I����W��_�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�d�e�f�m�G��I����V�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�l�G���Y���D��^�E��e�e�e�e�g�m�G��I����W��L����u�d�d�d�f�l�F��H����V��^�E��e�d�d�y�]�}�W��H����W��_�E��e�d�e�e�g�m�G��H���F�_�D��d�d�d�d�f�m�F��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�d�u�}�W���[����W��_�D��e�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��I����V��^�D��y�_�u�u�f�l�F��H����V��^�D��e�e�e�e�f�l�[�ԜY���W��_�D��e�e�d�d�f�m�G��I����W�d��U���d�d�d�d�f�l�G��I����V��^�E��d�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�F���Y���D��_�D��d�e�d�d�f�l�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�d�e�y�]�}�W��H����W��^�D��d�d�e�e�g�m�G��I���F�_�D��d�d�d�d�g�m�G��I����V��_�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�e�u�}�W���[����W��_�E��e�e�e�e�g�m�G��I����FǻN��D��d�d�d�d�g�l�F��I����V��^�D��y�_�u�u�f�l�F��H����W��^�D��e�e�e�e�f�l�[�ԜY���W��_�D��e�d�d�d�f�m�G��I����W�d��U���d�d�d�d�f�l�G��H����V��^�E��e�w�u�u�w��F��H����W��^�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�f�l�F��I����V��L����u�d�d�d�f�l�F��H����V��^�E��e�d�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�d�e�d�g�m�F��I����V��^�W���u�u�w�d�f�l�F��I����V��_�E��e�e�e�d�u�}�W���[����W��_�D��d�e�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��_�D��e�e�e�e�g�l�[�ԜY���W��_�D��d�e�d�e�f�m�G��I����V�d��U���d�d�d�d�f�m�F��I����V��^�E��d�w�u�u�w��F��H����V��^�D��d�e�e�e�g�m�F���Y���D��_�D��d�d�e�e�f�l�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��H���F�_�D��d�d�e�e�f�m�G��I����V��^�W���u�u�w�d�f�l�F��I����V��^�E��e�e�e�e�u�}�W���[����W��_�D��e�d�e�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��H����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��e�d�d�e�g�m�G��I����V�d��U���d�d�d�d�f�m�G��H����V��^�E��e�w�u�u�w��F��H����V��_�E��d�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�g�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��d�d�d�d�f�l�F��H���F�_�D��d�d�e�e�f�m�F��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��d�d�d�d�u�}�W���[����W��_�D��d�e�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��I����W��_�D��y�_�u�u�f�l�F��H����V��_�E��d�d�d�d�f�l�[�ԜY���W��_�D��d�e�d�e�f�l�F��H����V�d��U���d�d�d�d�f�m�F��I����W��_�D��d�w�u�u�w��F��H����V��^�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�e�e�g�m�F��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�e�y�]�}�W��H����W��_�D��e�e�d�d�f�l�F��I���F�_�D��d�d�e�d�f�l�G��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��d�d�d�d�u�}�W���[����W��_�D��d�e�e�e�f�l�F��H����FǻN��D��d�d�d�d�f�l�F��I����W��_�D��y�_�u�u�f�l�F��H����W��_�D��d�d�d�d�f�l�[�ԜY���W��_�D��d�d�e�d�g�l�F��H����W�d��U���d�d�d�d�f�m�F��H����W��_�D��e�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�G���Y���D��_�D��d�e�e�d�g�m�G��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�d�y�]�}�W��H����W��^�D��d�e�d�d�f�l�F��H���F�_�D��d�d�d�e�f�l�F��H����W��_�W���u�u�w�d�f�l�F��H����W��^�D��d�d�d�e�u�}�W���[����W��_�E��d�e�d�e�f�l�F��H����FǻN��D��d�d�d�d�g�l�G��H����W��_�D��y�_�u�u�f�l�F��H����W��_�D��d�d�d�d�f�m�[�ԜY���W��_�D��d�e�e�d�g�l�F��H����V�d��U���d�d�d�d�f�l�F��I����W��_�D��e�w�u�u�w��F��H����W��_�E��d�d�d�d�f�l�G���Y���D��_�D��d�e�e�d�g�m�G��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�e�y�]�}�W��H����W��^�E��e�e�d�d�f�l�F��I���F�_�D��d�d�d�d�g�l�F��H����W��_�W���u�u�w�d�f�l�F��H����W��^�D��d�d�d�e�u�}�W���[����W��_�E��d�d�d�e�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��I����W��_�D��y�_�u�u�f�l�F��H����V��^�D��d�d�d�d�f�m�[�ԜY���W��_�D��e�d�d�d�f�l�F��H����V�d��U���d�d�d�d�f�l�G��H����W��_�D��e�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�G���Y���D��_�D��d�d�d�d�f�l�F��H����W��L����u�d�d�d�f�l�F��H����V��_�D��d�d�e�y�]�}�W��H����W��_�D��e�d�d�d�f�l�F��I���F�_�D��d�d�d�d�g�m�G��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��d�d�d�e�u�}�W���[����W��_�D��e�e�e�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��H����W��_�D��y�_�u�u�f�l�F��H����V��_�E��d�d�d�d�f�l�[�ԜY���W��_�D��d�e�d�d�f�l�F��H����W�d��U���d�d�d�d�f�l�F��H����W��_�D��e�w�u�u�w��F��H����W��_�D��d�d�d�d�f�l�G���Y���D��_�D��d�d�d�d�g�l�G��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�d�d�y�]�}�W��I����V��^�E��e�d�d�d�f�l�F��H���F�^�E��e�e�e�e�g�l�G��H����W��_�W���u�u�w�e�g�m�G��I����V��^�D��d�d�d�e�u�}�W���[����V��^�E��d�e�d�d�f�l�F��H����FǻN��E��e�e�e�e�g�m�F��H����W��_�D��y�_�u�u�g�m�G��I����W��^�E��d�d�d�d�f�l�[�ԜY���V��^�E��e�e�e�d�g�l�F��H����W�d��U���e�e�e�e�g�m�G��H����W��_�D��e�w�u�u�w��G��I����V��_�E��e�d�d�d�f�l�G���Y���D��^�E��e�e�d�d�g�m�F��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�d�e�y�]�}�W��I����V��^�E��d�e�d�d�f�l�F��I���F�^�E��e�e�e�d�g�l�F��H����W��_�W���u�u�w�e�g�m�G��I����W��^�D��d�d�d�d�u�}�W���[����V��^�E��e�e�e�e�f�l�F��H����FǻN��E��e�e�e�e�g�m�G��I����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�f�m�[�ԜY���V��^�E��d�d�e�d�f�l�F��H����V�d��U���e�e�e�e�g�m�F��H����W��_�D��d�w�u�u�w��G��I����V��^�D��d�d�d�d�f�l�F���Y���D��^�E��e�e�d�e�f�m�F��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�d�e�y�]�}�W��I����V��^�E��e�e�d�d�f�l�F��H���F�^�E��e�e�e�d�g�l�G��H����W��_�W���u�u�w�e�g�m�G��I����V��^�D��d�d�d�d�u�}�W���[����V��^�E��e�d�d�e�f�l�F��H����FǻN��E��e�e�e�e�g�l�G��H����W��_�D��y�_�u�u�g�m�G��I����W��_�E��d�d�d�d�f�l�[�ԜY���V��^�E��d�d�e�d�g�l�F��H����W�d��U���e�e�e�e�g�m�F��I����W��_�D��d�w�u�u�w��G��I����V��_�E��e�d�d�d�f�l�F���Y���D��^�E��e�e�d�d�g�l�F��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�d�d�y�]�}�W��I����V��_�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�D��e�d�e�e�g�m�G��I����FǻN��E��e�e�e�e�f�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�G���Y���D��^�E��e�d�e�e�g�l�F��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��_�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�d�f�l�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�E��d�e�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�l�F��H����V��^�E��y�_�u�u�g�m�G��I����W��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�d�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�F��I����V��^�E��e�w�u�u�w��G��I����V��_�D��e�e�e�e�g�m�G���Y���D��^�E��e�e�d�e�g�m�F��I����V��L����u�e�e�e�g�m�G��H����W��^�E��e�e�d�y�]�}�W��I����V��^�D��d�d�e�e�g�m�G��H���F�^�E��e�e�e�d�g�l�F��I����V��^�W���u�u�w�e�g�m�G��I����W��_�E��e�e�e�e�u�}�W���[����V��^�E��d�d�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�l�F��I����V��^�E��y�_�u�u�g�m�G��I����W��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�e�d�e�f�m�G��I����W�d��U���e�e�e�e�g�m�F��I����V��^�E��e�w�u�u�w��G��I����V��_�D��d�e�e�e�g�m�G���Y���D��^�E��e�e�e�d�g�m�F��I����V��L����u�e�e�e�g�m�G��I����W��^�E��e�e�d�y�]�}�W��I����V��^�D��e�d�e�e�g�m�G��H���F�^�E��e�e�e�d�f�l�F��I����V��^�W���u�u�w�e�g�m�G��I����V��_�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�d�g�m�G��I����FǻN��E��e�e�e�e�g�m�F��I����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�e�d�d�f�m�G��I����W�d��U���e�e�e�e�g�m�F��H����V��^�E��e�w�u�u�w��G��I����V��^�D��d�e�e�e�g�m�G���Y���D��^�E��e�e�d�d�f�m�F��I����V��L����u�e�e�e�g�m�G��H����W��^�E��e�e�d�y�]�}�W��I����V��^�D��d�e�e�e�g�m�G��H���F�^�E��e�e�e�e�f�l�G��I����V��^�W���u�u�w�e�g�m�G��I����V��_�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�d�g�m�G��I����FǻN��E��e�e�e�e�g�l�F��I����V��^�E��y�_�u�u�g�m�G��I����W��_�D��e�e�e�e�g�l�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�G���Y���D��^�E��e�e�d�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����W��^�E��e�e�d�y�]�}�W��I����V��^�D��e�d�e�e�g�m�G��H���F�^�E��e�e�e�e�f�m�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�E��e�d�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��e�e�e�d�g�m�G��I����W�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�l�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�d�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��H���F�_�D��d�d�d�d�f�l�F��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�D��d�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��H����V��^�E��y�_�u�u�f�l�F��H����W��^�D��e�e�e�e�g�l�[�ԜY���W��_�D��d�d�d�e�g�m�G��I����W�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�E��d�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�f�l�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��e�e�d�y�]�}�W��H����W��_�E��d�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�D��e�d�e�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��I����V��^�E��y�_�u�u�f�l�F��H����W��^�D��e�e�e�e�g�l�[�ԜY���W��_�D��d�e�e�d�g�m�G��I����W�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�g�l�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�d�d�d�f�l�G��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�e�u�}�W���[����W��_�D��d�e�d�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�e�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�g�l�F��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�D��d�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�F��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�D��d�e�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��^�D��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�e�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�E��d�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�g�l�F��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�e�e�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�D��d�d�d�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�f�l�F��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�E��e�e�e�e�g�m�G��I���F�_�D��d�d�d�d�g�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�D��e�d�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��H����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�d�e�f�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��^�E��d�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�f�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�E��e�d�e�e�g�m�G��I���F�_�D��d�d�d�d�g�m�F��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�D��d�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��H����V��^�E��y�_�u�u�f�l�F��H����W��^�D��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��^�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�f�l�F��I����V��L����u�d�d�d�f�l�F��H����V��^�E��e�e�e�y�]�}�W��H����W��_�D��d�d�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�D��e�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��I����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�d�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�f�l�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��d�d�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�F��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�D��d�d�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��H����V��^�E��y�_�u�u�f�l�F��H����W��^�D��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�f�l�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��e�e�e�y�]�}�W��H����W��_�D��d�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�f�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��d�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�d�e�f�m�G��I����V�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��^�E��d�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��d�d�e�e�g�m�G��I���F�^�E��e�e�e�e�g�l�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�d�d�g�m�G��I����V�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��^�E��d�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W��E܍��V ��R����u�u�|�_�w�}�WϽ�����GF��X�����3��1�-�8�	����:����Z��P��O���u�u�x�i��*��������W��X������k�u�u�n�e�W���T����	��D�����;�0��'�?�.�6��s���l�T�����u��2�0�#�2��������A2��D#��D��<�!�2�'�m�}�W���T�ڧ�Z��D�����;�0��'�?�.�6��s���_��=N��U���z��2�0�#�2��������A2��D#��D�ߊu�u�_�u�8�.��������U+��X��U�����c�!�m�}�}���Y����p	��Q#�����k�u�u�_�w�}�G��I����V��^�E��e�e�e�e�g�m�G��U���F�^�E��e�e�e�e�g�m�G��I����V��^��U���u�w�e�e�g�m�G��I����V��^�E��e�e�e�w�w�}�W���I����V��^�E��e�e�e�e�g�m�G��I���9F�L�E��e�e�e�e�g�m�G��I����V��^�E���_�u�u�e�g�m�G��I����V��^�E��e�e�e�e�g�q�}���Y����V��^�E��e�e�e�e�g�m�G��I����J�N��W��e�e�e�e�g�m�G��I����V��^�E��w�u�u�u�u�m�G��I����V��^�E��e�e�e�e�g�m�U���Y���V��^�E��e�e�e�e�g�m�G��I����V��NךU���e�e�e�e�g�m�G��I����V��^�E��e�e�y�_�w�}�G��I����V��^�E��e�e�e�e�g�m�G��U���F�^�E��e�e�e�e�g�m�G��I����V��^��U���u�w�e�e�g�m�G��I����V��^�E��e�e�e�w�w�}�W���I����V��^�E��e�e�e�e�g�m�G��I���9F�L�E��e�e�e�e�g�m�G��I����V��^�E���_�u�u�e�g�m�G��I����V��^�E��e�e�e�e�g�q�}���Y����V��^�E��e�e�e�e�g�m�G��I����J�N��W��e�e�e�e�g�m�G��I����V��^�E��w�u�u�u�u�m�G��I����V��^�E��e�e�e�e�g�m�U���Y���V��^�E��e�e�e�e�g�m�G��I����V��NךU���e�e�e�e�g�m�G��I����V��^�E��e�e�y�_�w�}�G��I����V��^�E��e�e�e�e�g�m�G��U���F�^�E��e�e�e�e�g�m�G��I����V��^��U���u�w�e�e�g�m�G��I����V��^�E��e�e�e�w�w�}�W���I����V��^�E��e�e�e�e�g�m�G��I���9F�L�E��e�e�e�e�g�m�G��I����V��^�E���_�u�u�e�g�m�G��I����V��^�E��e�e�e�e�g�q�}���Y����V��^�E��e�e�e�e�g�m�G��I����J�N��W��e�e�e�e�g�m�G��I����V��^�E��w�u�u�u�u�m�G��I����V��^�E��e�e�e�e�g�m�U���Y���V��^�E��e�e�e�e�g�m�G��I����V��NךU���e�e�e�e�g�m�G��I����V��^�E��e�e�y�_�w�}�G��I����V��^�E��e�e�e�e�g�m�G��U���F�^�E��e�e�e�e�g�m�G��I����V��^��U���u�w�e�e�g�m�G��I����V��^�E��e�e�e�w�w�}�W���I����V��^�E��e�e�e�e�g�m�G��I���9F�L�E��e�e�e�e�g�m�G��I����V��^�E���_�u�u�e�g�m�G��I����V��^�E��e�e�e�e�g�q�}���Y����V��^�E��e�e�e�e�g�m�G��I����J�N��W��e�e�e�e�g�m�G��I����V��^�E��w�u�u�u�u�m�G��I����V��^�E��e�e�e�e�g�m�U���Y���V��^�E��e�e�e�e�g�m�G��I����V��NךU���e�e�e�e�g�m�G��I����V��^�E��e�e�y�_�w�}�G��I����V��^�E��e�e�e�e�g�m�G��U���F�^�E��e�e�e�e�g�m�G��I����V��^��U���u�w�e�e�g�m�G��I����V��^�E��e�e�e�w�w�}�W���I����W��^�D��e�e�e�d�f�l�F��H���9F�L�E��d�d�d�e�g�l�F��I����W��^�E���_�u�u�e�g�m�F��H����V��^�D��d�d�e�d�f�q�}���Y����V��_�E��d�d�d�d�f�l�F��H����J�N��W��e�e�d�d�g�l�F��H����W��_�D��w�u�u�u�u�m�G��H����V��^�D��d�d�d�d�g�l�U���Y���V��^�D��d�e�e�d�f�m�F��H����W��NךU���e�e�e�d�f�m�F��H����V��_�D��e�d�y�_�w�}�G��I����V��_�E��d�d�d�d�f�l�G��U���F�^�E��d�e�d�e�g�l�F��I����V��^��U���u�w�e�e�g�l�F��H����W��^�E��e�d�d�w�w�}�W���I����W��^�D��d�e�d�e�g�m�G��H���9F�L�E��d�d�e�e�f�m�F��I����V��_�E���_�u�u�e�g�m�F��I����V��_�E��e�e�e�e�g�q�}���Y����V��_�D��d�d�e�d�g�m�G��I����J�N��W��e�e�d�e�f�l�F��I����V��^�E��w�u�u�u�u�m�G��H����V��_�E��e�e�e�d�f�l�U���Y���V��^�D��d�e�e�e�g�l�G��I����W��NךU���e�e�e�d�f�m�F��H����V��^�D��e�d�y�_�w�}�G��I����V��^�D��e�e�e�e�f�l�G��U���F�^�E��e�e�e�d�g�m�G��I����W��_��U���u�w�e�e�g�l�F��H����V��^�E��d�e�d�w�w�}�W���I����W��^�D��e�e�e�e�g�m�F��H���9F�L�E��d�e�d�e�g�l�F��H����V��^�D���_�u�u�e�g�m�F��I����W��^�E��e�d�d�e�f�q�}���Y����V��^�E��d�d�e�d�g�m�G��I����J�N��W��e�e�d�e�f�m�G��I����V��^�D��w�u�u�u�u�m�G��H����W��^�D��e�e�d�e�g�l�U���Y���V��^�E��d�d�e�d�f�l�G��H����W��NךU���e�e�e�d�f�l�G��I����V��^�E��e�d�y�_�w�}�G��I����W��^�E��d�e�e�e�g�m�G��U���F�^�E��d�e�e�d�g�m�F��I����W��^��U���u�w�e�e�g�m�G��H����W��^�E��d�d�e�w�w�}�W���I����V��_�E��d�e�d�e�g�l�F��H���9F�L�E��d�d�e�e�f�l�F��H����W��^�E���_�u�u�e�g�m�F��H����V��^�E��e�d�e�d�g�q�}���Y����V��^�E��d�e�d�d�g�m�G��H����J�N��W��e�e�e�e�f�l�G��I����V��_�D��w�u�u�u�u�m�G��I����V��^�E��e�e�d�d�g�m�U���Y���V��^�D��d�d�d�d�g�l�G��H����W��NךU���e�e�e�e�f�m�F��I����W��^�D��d�e�y�_�w�}�G��I����W��_�D��d�e�e�e�f�l�G��U���F�^�E��e�e�e�e�f�m�G��I����W��^��U���u�w�e�e�g�l�G��I����W��^�E��d�d�e�w�w�}�W���I����W��^�E��d�d�e�e�g�m�G��H���9F�L�E��e�e�d�d�f�l�F��I����V��_�E���_�u�u�e�g�m�G��I����V��_�E��d�e�e�d�g�q�}���Y����V��_�D��e�d�e�d�g�m�F��H����J�N��W��e�e�e�d�f�m�F��I����V��^�E��w�u�u�u�u�m�G��I����W��_�E��e�e�e�e�f�m�U���Y���V��^�D��e�d�d�e�f�m�G��I����V��NךU���e�e�e�e�g�l�F��H����W��^�E��e�d�y�_�w�}�G��I����V��_�E��e�e�e�d�g�m�F��U���F�^�E��e�e�d�d�f�m�G��I����V��_��U���u�w�e�e�g�m�G��I����V��^�E��d�d�d�w�w�}�W���H����W��_�D��d�d�e�e�g�m�F��I���9F�L�D��d�d�d�e�g�l�G��H����V��_�D���_�u�u�d�f�l�F��I����V��_�E��d�e�d�e�f�q�}���Y����W��^�E��e�e�e�e�g�m�F��H����J�N��W��d�d�d�d�g�m�F��I����V��^�E��w�u�u�u�u�l�F��H����V��^�E��e�e�e�d�g�m�U���Y���W��_�D��e�e�e�e�f�l�G��I����W��NךU���d�d�d�d�f�m�F��H����V��^�E��d�e�y�_�w�}�F��H����W��_�D��e�e�e�d�g�l�F��U���F�_�D��e�e�e�e�g�m�G��I����W��^��U���u�w�d�d�f�m�F��I����V��^�E��d�e�d�w�w�}�W���H����V��_�D��d�d�e�e�g�m�F��I���9F�L�D��d�e�e�d�g�m�F��H����V��^�E���_�u�u�d�f�l�G��H����W��_�E��d�e�d�e�g�q�}���Y����W��_�D��d�d�e�d�g�m�F��H����J�N��W��d�d�d�e�f�m�F��I����V��^�D��w�u�u�u�u�l�F��H����W��_�E��e�e�e�d�f�m�U���Y���W��_�E��d�d�e�d�f�l�G��I����W��NךU���d�d�d�e�g�l�F��I����V��^�E��d�d�y�_�w�}�F��H����V��^�D��d�e�e�d�g�m�G��U���F�_�D��d�e�e�d�f�l�F��I����V��^��U���u�w�d�d�f�m�G��H����W��^�E��e�d�e�w�w�}�W���H����V��_�D��e�e�e�e�g�m�G��H���9F�L�D��e�e�d�d�g�m�F��H����V��^�D���_�u�u�d�f�l�G��I����V��_�E��d�e�e�d�g�q�}���Y����W��^�D��e�d�e�e�g�m�F��I����J�N��W��d�d�e�e�f�l�F��H����V��^�E��w�u�u�u�u�l�F��H����W��_�E��e�e�d�d�f�m�U���Y���W��^�D��e�d�e�d�f�m�G��H����W��NךU���d�d�d�d�f�l�F��I����W��^�D��e�d�y�_�w�}�F��H����V��^�E��d�e�e�e�f�m�G��U���F�_�E��d�d�d�d�g�l�G��I����V��_��U���u�w�d�d�g�l�F��H����V��^�E��e�d�e�w�w�}�W���H����W��^�E��e�e�e�e�g�l�G��I���9F�L�D��d�e�d�e�g�m�G��H����W��_�E���_�u�u�d�f�l�F��I����W��^�E��e�d�e�d�g�q�}���Y����W��^�E��e�d�d�e�g�m�G��H����J�N��W��d�e�e�d�g�m�F��H����V��^�E��w�u�u�u�u�l�F��I����W��^�D��e�e�d�d�f�l�U���Y���W��^�D��e�e�d�d�g�l�G��H����V��NךU���d�d�d�d�f�l�F��H����V��^�E��d�d�y�_�w�}�F��H����V��^�E��d�e�e�e�g�m�F��U���F�_�E��e�e�e�d�g�m�F��I����V��^��U���u�w�d�d�g�m�F��H����W��^�E��d�d�d�w�w�}�W���H����V��^�D��d�d�e�e�g�m�F��H���9F�L�D��d�e�d�e�g�l�G��H����V��^�D���_�u�u�d�f�l�F��I����W��_�E��e�d�d�e�g�q�}���Y����W��^�E��e�e�e�d�g�m�G��I����J�N��W��d�e�e�d�g�l�G��I����V��_�E��w�u�u�u�u�l�F��I����W��^�E��e�e�e�d�f�m�U���Y���W��^�E��e�d�e�e�g�m�G��I����W��NךU���d�d�d�d�g�l�G��I����W��^�E��e�e�y�_�w�}�F��H����W��^�D��e�e�e�e�g�l�F��U���F�_�E��e�e�d�e�f�m�F��I����V��_��U���u�w�d�d�g�m�G��H����W��_�D��d�d�d�w�w�}�W���H����V��_�E��e�e�e�d�f�l�F��H���9F�L�D��d�e�d�e�f�l�F��I����W��^�D���_�u�u�d�f�l�F��H����W��_�D��d�d�d�e�g�q�}���Y����W��^�D��e�d�d�d�f�l�F��I����J�N��W��d�e�e�d�g�l�G��H����W��_�E��w�u�u�u�u�l�F��I����W��_�E��d�d�d�d�g�l�U���Y���W��^�E��d�d�d�e�g�m�F��H����V��NךU���d�d�d�d�g�l�G��I����W��_�E��d�d�y�_�w�}�F��H����W��^�E��e�d�d�d�g�l�G��U���F�_�E��e�e�d�e�g�l�F��H����V��^��U���u�w�d�d�g�m�G��H����V��_�D��d�d�e�w�w�}�W���H����V��^�E��e�e�d�d�f�m�F��H���9F�L�D��d�d�d�d�g�m�F��I����V��_�D���_�u�u�d�f�l�F��I����V��^�D��d�d�d�e�f�q�}���Y����W��_�E��d�d�e�e�f�l�F��I����J�N��W��d�e�d�e�g�m�G��I����W��^�D��w�u�u�u�u�l�F��H����W��^�D��d�d�e�d�f�l�U���Y���W��^�E��e�d�d�d�g�l�F��I����W��NךU���d�d�d�d�g�m�G��I����W��_�E��d�e�y�_�w�}�F��H����W��_�D��e�d�d�d�g�m�G��U���F�_�E��e�d�e�d�f�m�G��H����W��_��U���u�w�d�d�g�l�G��H����W��_�D��d�e�e�w�w�}�W���H����W��_�E��d�e�e�d�f�l�F��I���9F�L�D��d�d�d�d�g�l�F��I����W��_�D���_�u�u�d�f�l�G��H����V��_�D��e�d�d�e�f�q�}���Y����W��^�E��d�d�e�d�f�l�G��I����J�N��W��d�d�e�d�f�m�F��I����W��^�D��w�u�u�u�u�l�F��I����V��_�D��d�d�d�d�g�l�U���Y���W��_�D��e�d�e�d�f�m�F��H����V��NךU���d�d�d�e�f�l�G��I����W��_�E��d�d�y�_�w�}�F��H����V��_�E��d�d�d�e�g�l�F��U���F�_�D��d�e�d�d�f�l�G��H����V��_��U���u�w�d�d�f�l�F��H����W��_�D��e�e�e�w�w�}�W���H����W��^�D��e�d�d�d�f�m�F��H���9F�L�D��e�d�e�d�f�l�G��I����V��^�D���_�u�u�d�f�l�F��I����V��^�D��e�d�e�e�f�q�}���Y����W��^�E��e�e�e�e�f�l�G��I����J�N��W��d�d�e�d�f�m�G��I����W��_�D��w�u�u�u�u�l�F��I����W��_�D��d�d�e�e�g�m�U���Y���W��_�D��e�d�e�d�g�m�F��I����W��NךU���d�d�d�d�g�m�F��I����V��_�D��e�e�y�_�w�}�F��H����V��^�D��e�d�d�e�f�m�G��U���F�_�D��e�e�d�d�f�m�F��H����W��_��U���u�w�d�d�f�l�F��H����W��_�D��d�d�e�w�w�}�W���I����V��^�E��e�e�e�d�f�m�F��H���9F�L�E��e�e�d�d�f�m�F��I����V��_�D���_�u�u�e�g�m�G��H����W��^�D��e�e�e�e�f�q�}���Y����V��_�E��d�d�e�e�f�l�G��I����J�N��W��e�e�e�d�g�m�F��H����W��^�E��w�u�u�u�u�m�G��H����W��^�E��d�d�e�d�g�l�U���Y���V��^�E��e�d�e�d�f�m�F��I����V��NךU���e�e�e�e�f�m�F��I����V��_�E��d�e�y�_�w�}�G��I����V��_�D��d�d�d�e�g�l�F��U���F�^�E��e�d�e�e�g�l�G��H����W��^��U���u�w�e�e�g�m�F��H����W��_�D��e�d�e�w�w�}�W���I����V��_�E��d�d�e�d�f�m�G��I���9F�L�E��d�d�e�d�g�l�G��H����V��_�D���_�u�u�e�g�m�F��I����W��^�D��e�e�d�d�g�q�}���Y����V��^�E��d�e�d�d�f�l�G��I����J�N��W��e�e�d�e�g�m�F��H����W��^�E��w�u�u�u�u�m�G��H����W��_�D��d�d�e�d�g�m�U���Y���V��^�D��e�d�d�e�g�m�F��I����V��NךU���e�e�e�e�g�l�G��I����W��_�E��d�e�y�_�w�}�G��I����W��^�D��e�d�d�e�g�l�G��U���F�^�D��e�e�d�d�f�m�F��H����W��_��U���u�w�e�e�f�m�F��H����V��_�D��d�d�d�w�w�}�W���I����W��_�D��e�e�e�d�f�m�G��I���9F�L�E��e�e�e�d�g�l�G��I����V��^�E���_�u�u�e�g�m�G��I����V��_�D��e�d�e�d�g�q�}���Y����V��_�D��d�d�d�e�f�l�G��H����J�N��W��e�d�d�d�g�l�G��H����W��_�D��w�u�u�u�u�m�G��I����V��^�E��d�d�e�d�g�l�U���Y���V��_�E��e�e�e�d�f�l�F��I����V��NךU���e�e�e�d�f�m�G��H����V��_�D��d�d�y�_�w�}�G��I����W��^�D��d�d�d�e�f�l�F��U���F�^�D��d�e�d�e�f�m�G��H����V��_��U���u�w�e�e�f�l�G��I����W��_�D��e�e�d�w�w�}�W���I����W��_�D��d�e�e�d�f�l�G��H���9F�L�E��d�e�d�d�g�m�F��H����W��_�E���_�u�u�e�g�m�F��I����W��_�D��e�e�d�d�g�q�}���Y����V��_�D��e�d�e�d�f�l�G��I����J�N��W��e�d�d�d�g�m�G��I����W��_�D��w�u�u�u�u�m�G��I����W��^�E��d�d�d�e�f�m�U���Y���V��^�E��e�d�d�e�g�m�F��H����W��NךU���e�e�d�e�g�m�F��H����V��_�D��e�e�y�_�w�}�G��H����W��_�D��d�d�d�d�g�m�F��U���F�^�E��e�e�d�d�f�l�G��H����W��_��U���u�w�e�e�g�m�G��I����V��_�D��d�e�e�w�w�}�W���I����V��_�D��e�e�e�d�f�m�F��I���9F�L�E��e�d�e�e�g�l�G��I����V��^�E���_�u�u�e�g�l�G��H����V��^�D��d�d�d�d�g�q�}���Y����W��_�D��e�e�d�e�f�l�F��I����J�N��W��e�e�d�e�g�l�G��I����W��_�E��w�u�u�u�u�m�G��H����V��^�E��d�d�d�e�g�l�U���Y���V��^�E��d�e�e�e�g�m�F��H����V��NךU���e�e�d�e�g�l�G��H����V��_�E��e�e�y�_�w�}�G��H����W��_�D��e�d�d�d�g�l�F��U���F�^�E��d�e�e�d�f�m�F��H����V��_��U���u�w�e�e�g�l�F��H����V��_�D��d�e�e�w�w�}�W���I����W��^�D��e�e�e�d�f�l�F��I���9F�L�E��e�e�e�e�g�l�F��I����V��^�D���_�u�u�e�g�l�G��I����W��_�E��e�e�d�e�g�q�}���Y����W��^�D��e�d�e�d�g�m�G��I����J�N��W��e�e�d�e�f�l�G��I����V��_�E��w�u�u�u�u�m�G��H����V��^�D��e�e�e�e�g�m�U���Y���V��^�E��d�e�e�d�f�m�G��I����V��NךU���e�e�d�e�g�m�F��H����W��^�D��d�e�y�_�w�}�G��H����W��_�E��d�e�e�e�g�l�G��U���F�^�E��d�e�d�d�g�l�F��I����V��^��U���u�w�e�e�g�m�F��I����V��^�E��d�d�e�w�w�}�W���I����V��_�D��d�d�d�e�g�l�G��I���9F�L�E��e�d�e�d�f�m�F��H����W��^�E���_�u�u�e�g�l�G��H����W��_�E��e�d�d�d�f�q�}���Y����W��^�D��e�d�e�d�g�m�F��I����J�N��W��e�e�e�e�f�l�F��H����V��^�D��w�u�u�u�u�m�G��I����V��^�D��e�e�e�d�g�m�U���Y���V��_�D��d�e�d�e�f�l�G��I����V��NךU���e�e�e�d�f�l�F��H����V��^�D��e�e�y�_�w�}�G��I����V��^�E��e�e�e�d�f�m�F��U���F�^�D��d�e�e�e�g�l�G��I����W��_��U���u�w�e�e�f�l�G��H����W��^�E��e�e�d�w�w�}�W���I����V��_�E��d�d�e�e�g�l�F��H���9F�L�E��d�d�e�e�g�l�G��H����W��_�D���_�u�u�e�g�m�F��I����V��^�E��d�d�e�d�g�q�}���Y����V��^�E��e�e�e�e�g�m�F��H����J�N��W��e�d�e�e�g�l�G��H����V��_�E��w�u�u�u�u�m�G��H����W��_�E��e�d�e�e�g�l�U���Y���V��_�D��d�d�d�e�g�l�G��I����V��NךU���e�e�e�e�g�m�G��I����V��_�E��d�d�y�_�w�}�G��I����V��^�D��e�e�e�e�g�l�F��U���F�^�D��e�d�d�d�f�l�F��I����V��_��U���u�w�e�e�f�m�F��H����V��^�D��e�e�d�w�w�}�W���I����V��_�D��d�d�d�e�f�m�F��H���9F�L�E��d�d�e�e�g�l�F��I����V��^�E���_�u�u�e�g�m�F��I����V��^�E��e�e�e�d�f�q�}���Y����V��^�E��d�e�d�e�g�m�G��H����J�N��W��e�e�e�d�f�m�F��H����V��^�E��w�u�u�u�u�m�G��I����V��_�D��e�d�d�d�g�m�U���Y���V��^�E��d�d�d�d�f�l�G��H����V��NךU���e�e�e�e�f�m�G��H����V��_�D��e�d�y�_�w�}�G��I����W��^�E��d�e�e�e�f�l�F��U���F�^�E��e�d�d�e�g�m�F��I����V��_��U���u�w�e�e�g�m�G��H����W��^�D��d�d�d�w�w�}�W���I����V��_�D��d�d�d�e�f�l�F��H���9F�L�E��e�e�e�e�g�m�G��I����W��_�D���_�u�u�d�f�l�F��I����W��^�E��d�e�e�e�g�q�}���Y����W��^�D��e�d�e�e�g�m�F��H����J�N��W��d�d�e�d�f�m�F��H����V��^�D��w�u�u�u�u�l�F��I����W��_�D��e�d�e�e�f�l�U���Y���W��_�E��e�e�e�d�g�m�G��I����W��NךU���d�d�d�e�f�l�F��H����W��_�E��e�d�y�_�w�}�F��H����V��^�E��e�e�e�d�g�l�G��U���F�_�D��d�d�d�d�g�m�F��I����W��_��U���u�w�d�d�f�m�F��I����V��^�D��d�d�e�w�w�}�W���H����V��_�E��e�d�e�e�f�m�F��H���9F�L�D��d�d�d�d�g�m�F��I����V��_�D���_�u�u�d�f�l�F��I����V��_�E��d�e�d�d�g�q�}���Y����W��_�D��d�e�e�d�g�m�F��H����J�N��W��d�e�e�d�f�m�F��I����V��^�D��w�u�u�u�u�l�F��I����V��_�E��e�d�e�d�f�m�U���Y���W��^�D��e�d�d�d�f�l�G��I����W��NךU���d�d�d�e�g�l�F��H����W��_�E��e�e�y�_�w�}�F��H����V��^�D��d�e�e�d�g�l�F��U���F�_�E��d�e�d�d�f�m�F��I����W��^��U���u�w�d�d�g�m�G��I����W��^�D��d�d�d�w�w�}�W���H����W��^�E��e�d�e�e�f�m�F��I���9F�L�D��d�e�e�e�g�l�G��I����V��_�E���_�u�u�d�f�m�F��I����V��_�E��d�e�d�d�g�q�}���Y����V��^�D��d�d�d�e�g�m�F��I����J�N��W��d�d�e�e�f�l�F��I����V��^�E��w�u�u�u�u�l�F��H����W��_�D��e�d�d�d�f�m�U���Y���W��_�E��e�e�e�e�f�m�G��H����W��NךU���d�d�e�e�g�m�G��H����W��_�D��e�e�y�_�w�}�F��I����W��^�D��e�e�e�e�f�l�F��U���F�_�D��d�d�e�e�f�l�G��I����V��_��U���u�w�d�d�g�l�F��I����V��^�D��d�d�e�w�w�}�W���H����W��^�E��d�d�e�e�f�l�F��I���9F�L�D��d�e�e�e�g�m�G��I����W��_�D���_�u�u�d�f�m�F��I����V��^�E��e�e�e�d�f�q�}���Y����V��_�D��d�d�d�e�g�m�G��H����J�N��W��d�e�e�d�g�l�F��I����V��_�E��w�u�u�u�u�l�F��I����V��_�D��e�d�e�e�f�l�U���Y���W��^�D��e�e�e�e�g�m�G��I����W��NךU���d�d�e�e�f�m�F��I����W��_�E��d�d�y�_�w�}�F��I����V��^�E��d�e�e�e�g�m�F��U���F�_�E��e�e�d�e�g�l�F��I����W��^��U���u�w�d�d�g�m�F��I����W��^�E��d�e�e�w�w�}�W���H����V��_�E��d�e�d�e�g�l�G��H���9F�L�D��e�e�d�e�f�l�F��I����W��_�E���_�u�u�d�f�m�G��H����V��_�E��d�e�d�d�g�q�}���Y����V��^�E��e�e�d�d�g�m�F��H����J�N��W��e�d�d�d�f�l�G��H����V��_�D��w�u�u�u�u�l�G��H����W��_�E��e�e�e�e�g�m�U���Y���W��_�D��d�e�d�e�g�l�G��I����V��NךU���d�d�d�d�g�l�F��H����W��^�E��d�d�y�_�w�}�F��H����V��_�D��d�e�e�e�f�m�G��U���F�_�D��e�d�e�e�g�l�G��I����V��_��U���u�w�d�e�f�l�G��H����W��^�E��d�d�d�w�w�}�W���H����W��^�E��e�d�e�e�g�l�G��I���9F�L�D��d�d�d�d�f�m�F��I����V��_�D���_�u�u�d�f�l�F��H����V��_�E��e�d�e�d�f�q�}���Y����W��_�D��d�e�d�d�g�m�G��I����J�N��W��e�d�e�d�f�m�F��H����V��^�E��w�u�u�u�u�l�G��I����W��^�D��d�d�d�e�f�l�U���Y���W��_�D��d�d�e�e�f�m�F��H����V��NךU���d�d�d�d�g�m�F��I����W��_�E��d�d�y�_�w�}�F��H����V��^�D��e�d�d�d�f�l�G��U���F�_�D��e�d�e�d�g�m�F��H����V��^��U���u�w�d�e�f�l�F��H����V��_�D��d�d�e�w�w�}�W���H����W��^�E��e�d�d�d�f�m�G��H���9F�L�D��d�d�e�e�f�m�G��H����W��_�E���_�u�u�d�f�l�F��H����W��^�D��e�e�d�d�f�q�}���Y����W��_�E��d�d�e�d�f�l�G��I����J�N��W��d�e�e�e�f�l�F��I����W��_�E��w�u�u�u�u�l�F��I����W��^�D��d�d�e�e�g�m�U���Y���W��^�D��e�d�e�e�g�l�F��I����V��NךU���d�d�e�e�f�m�G��I����V��^�D��e�e�y�_�w�}�F��I����V��_�E��d�d�d�d�f�m�G��U���F�_�E��d�e�d�d�f�m�G��H����W��_��U���u�w�d�d�g�l�G��I����V��_�E��d�e�d�w�w�}�W���H����V��^�D��d�d�e�d�g�m�G��H���9F�L�D��d�e�d�d�g�l�F��H����V��^�D���_�u�u�d�f�m�F��I����V��_�D��e�d�d�d�f�q�}���Y����V��^�E��d�d�d�e�f�l�G��H����J�N��W��d�e�d�e�f�m�G��H����W��^�D��w�u�u�u�u�l�F��I����V��_�D��d�e�d�e�g�l�U���Y���W��_�E��d�d�e�d�g�m�F��I����V��NךU���d�d�e�e�f�l�F��I����V��^�E��e�d�y�_�w�}�F��I����W��^�E��e�d�d�e�g�m�G��U���F�_�D��d�d�d�e�g�m�F��I����V��^��U���u�w�d�d�f�m�G��H����W��_�D��d�e�d�w�w�}�W���H����W��_�D��e�d�d�d�f�l�G��H���9F�L�D��d�d�d�e�f�m�G��I����V��_�E���_�u�u�d�f�l�G��H����V��_�D��d�d�e�e�g�q�}���Y����W��_�D��d�d�e�e�f�m�F��H����J�N��W��d�e�d�d�f�l�F��H����V��_�E��w�u�u�u�u�l�F��I����V��^�D��d�d�d�e�f�l�U���Y���W��^�D��d�d�e�e�g�l�F��H����V��NךU���d�d�d�d�g�l�F��I����W��_�D��d�d�y�_�w�}�F��H����W��_�D��d�d�e�e�f�l�G��U���F�_�D��d�e�d�d�f�m�G��I����W��_��U���u�w�d�d�f�l�G��I����V��_�D��e�e�e�w�w�}�W���H����V��^�E��e�d�e�d�g�l�F��I���9F�L�D��d�e�d�e�g�l�G��I����W��_�D���_�u�u�e�g�m�G��I����V��^�D��d�e�e�d�g�q�}���Y����V��_�E��d�e�e�d�f�m�F��I����J�N��W��e�e�d�e�g�m�F��I����V��_�E��w�u�u�u�u�m�G��I����V��^�D��d�e�e�e�g�m�U���Y���V��^�E��e�d�d�d�g�l�F��I����V��NךU���e�e�e�e�g�l�G��H����V��^�E��e�d�y�_�w�}�G��I����V��_�D��d�d�e�e�f�m�G��U���F�^�D��e�e�e�d�f�m�G��I����V��_��U���u�w�e�e�f�m�F��H����W��_�E��d�e�d�w�w�}�W���I����W��_�D��e�d�e�d�g�l�G��H���9F�L�E��e�d�e�d�g�l�F��I����V��_�D���_�u�u�e�g�l�G��I����V��^�D��e�d�d�d�g�q�}���Y����W��_�D��d�d�d�d�f�m�G��H����J�N��W��e�e�d�e�f�l�F��I����V��^�E��w�u�u�u�u�m�G��I����W��_�E��d�e�e�e�f�l�U���Y���V��_�D��d�e�e�d�g�m�G��H����W��NךU���e�e�d�d�f�l�F��H����V��_�D��d�e�y�_�w�}�G��H����V��_�E��e�d�d�d�f�m�F��U���F�^�E��d�e�d�d�f�l�F��H����W��_��U���u�w�e�d�g�l�F��I����V��_�D��d�e�e�w�w�}�W���I����V��^�D��d�d�e�e�f�l�G��H���9F�L�E��d�d�d�d�g�m�G��H����V��_�D���_�u�u�e�g�m�G��I����V��_�D��d�d�e�d�f�q�}���Y����V��^�D��e�e�d�e�f�l�F��H����J�N��W��d�d�d�e�f�l�G��H����W��_�E��w�u�u�u�u�m�F��I����W��^�D��e�d�e�e�g�m�U���Y���V��^�E��e�e�e�d�g�m�G��I����V��NךU���e�e�d�d�g�l�F��I����V��_�E��d�e�y�_�w�}�G��H����V��_�D��d�d�d�d�g�m�F��U���F�^�D��e�d�d�d�f�m�G��H����W��_��U���u�w�e�d�f�l�F��H����V��_�D��e�e�d�w�w�}�W���I����V��_�D��d�d�d�e�f�m�G��I���9F�L�D��e�e�e�e�g�l�F��H����V��_�E���_�u�u�e�f�m�G��H����W��^�D��d�e�e�e�f�q�}���Y����V��^�E��e�d�d�d�f�l�F��I����J�N��W��e�e�d�d�g�l�G��I����W��^�E��w�u�u�u�u�m�G��I����W��^�E��e�d�e�e�g�l�U���Y���V��_�D��d�e�e�e�g�l�G��I����V��NךU���e�d�e�d�f�m�F��I����V��_�E��d�e�y�_�w�}�G��I����W��^�D��d�d�d�d�g�l�G��U���F�_�E��e�e�d�d�g�m�G��H����W��^��U���u�w�e�e�g�m�G��I����V��_�D��e�d�e�w�w�}�W���I����W��_�E��d�e�d�e�f�m�F��I���9F�L�D��e�e�e�e�f�l�G��I����V��_�D���_�u�u�e�f�l�G��H����V��_�D��d�e�d�e�f�q�}���Y����W��_�E��d�d�e�e�f�l�F��I����J�N��W��e�d�d�e�f�l�F��H����W��_�E��w�u�u�u�u�m�F��I����V��_�E��e�d�e�d�g�m�U���Y���V��^�D��e�d�e�e�g�l�G��I����V��NךU���e�d�e�d�f�m�G��I����W��_�E��e�d�y�_�w�}�G��I����W��^�E��d�d�d�d�g�l�F��U���F�_�D��d�e�e�d�f�l�F��H����V��_��U���u�w�e�d�f�l�F��H����V��_�D��d�d�e�w�w�}�W���I����V��_�D��d�d�d�e�f�l�G��H���9F�L�D��d�d�d�d�g�m�G��I����W��_�D���_�u�u�e�f�l�G��H����V��^�D��e�e�e�e�f�q�}���Y����W��_�D��d�e�d�d�f�m�G��H����J�N��W��d�e�e�d�f�m�F��H����V��^�E��w�u�u�u�u�m�F��H����V��_�D��d�e�e�e�g�m�U���Y���V��_�D��d�d�e�e�g�l�F��I����W��NךU���e�d�d�e�f�m�F��H����W��^�E��d�e�y�_�w�}�G��H����W��^�D��d�d�e�e�g�m�G��U���F�_�D��e�d�e�d�g�m�F��I����V��_��U���u�w�d�e�g�m�F��H����V��_�E��d�d�e�w�w�}�W���H����W��_�D��e�d�d�d�g�m�G��H���9F�L�E��d�e�d�e�g�m�F��H����V��^�D���_�u�u�e�g�m�F��I����V��^�D��d�d�d�d�f�q�}���Y����V��_�D��e�e�d�e�f�m�F��H����J�N��W��e�d�e�e�g�l�G��H����V��^�E��w�u�u�u�u�l�G��H����W��_�E��d�e�d�e�f�l�U���Y���W��_�E��d�d�d�e�f�l�F��H����W��NךU���e�e�e�d�f�l�F��H����W��_�E��d�d�y�_�w�}�G��I����W��_�E��d�d�e�e�f�m�F��U���F�^�E��d�d�e�d�f�l�F��I����W��^��U���u�w�d�e�g�l�G��I����W��_�D��e�d�d�w�w�}�W���H����W��^�D��d�d�e�d�f�l�G��H���9F�L�E��d�e�e�e�f�l�F��H����W��_�D���_�u�u�e�g�l�F��H����W��_�D��d�e�e�d�f�q�}���Y����W��^�D��e�e�e�e�f�m�F��H����J�N��W��e�d�e�e�g�l�F��I����V��^�E��w�u�u�u�u�l�G��I����V��_�E��d�d�d�d�g�l�U���Y���W��_�E��e�d�e�d�f�l�F��H����V��NךU���e�e�d�e�f�m�G��I����V��^�E��e�e�y�_�w�}�G��H����V��_�D��e�d�d�e�f�m�F��U���F�^�D��d�d�d�e�f�l�G��H����W��_��U���u�w�d�e�f�m�F��I����V��_�E��d�e�d�w�w�}�W���H����W��^�D��d�e�e�d�g�l�F��H���9F�L�E��d�d�d�e�g�m�F��I����V��_�D���_�u�u�e�g�l�F��H����V��^�D��d�d�d�e�f�q�}���Y����V��^�E��d�d�e�d�f�l�F��I����J�N��W��d�e�e�e�g�l�F��I����W��^�D��w�u�u�u�u�l�F��I����W��^�D��d�e�d�d�g�l�U���Y���W��^�E��d�d�d�e�f�l�F��I����V��NךU���e�e�e�e�g�l�F��H����V��_�D��d�d�y�_�w�}�G��I����W��_�D��e�d�d�e�g�l�F��U���F�^�E��e�d�e�e�g�l�G��H����V��^��U���u�w�d�d�g�l�G��I����W��_�D��e�e�e�w�w�}�W���H����W��^�D��e�e�e�d�f�m�F��I���9F�L�E��e�d�e�d�f�m�F��I����V��^�E���_�u�u�e�g�m�G��H����W��_�D��d�e�e�d�g�q�}���Y����V��_�E��d�d�e�d�f�l�F��I����J�N��W��d�e�d�d�g�l�F��I����V��^�D��w�u�u�u�u�l�F��H����V��_�E��e�e�e�e�g�m�U���Y���W��^�D��d�d�e�e�g�m�G��H����V��NךU���e�e�e�e�f�l�G��H����W��^�D��e�d�y�_�w�}�G��I����V��_�E��e�e�e�e�f�l�G��U���F�^�E��d�e�e�d�f�m�G��I����W��^��U���u�w�d�d�g�l�G��H����W��^�E��d�d�d�w�w�}�W���H����W��^�D��e�d�d�e�g�l�F��I���9F�L�E��e�d�e�d�f�l�F��H����W��_�E���_�u�u�e�g�m�G��I����W��_�E��e�e�e�d�g�q�}���Y����V��^�E��d�d�e�d�g�m�G��I����J�N��W��e�d�d�d�f�l�G��I����V��_�D��w�u�u�u�u�l�G��H����V��^�E��e�d�d�d�f�l�U���Y���W��_�E��e�d�d�d�g�m�G��H����V��NךU���e�e�d�d�f�l�G��H����V��_�E��e�d�y�_�w�}�G��H����W��_�D��e�e�e�d�f�m�F��U���F�^�D��e�e�d�e�f�m�G��I����V��_��U���u�w�d�e�f�l�G��I����V��^�D��d�e�e�w�w�}�W���H����W��_�D��d�d�d�e�f�l�F��H���9F�L�E��e�d�e�e�g�m�F��I����V��_�E���_�u�u�e�g�l�G��I����V��^�E��e�d�e�e�f�q�}���Y����W��^�D��e�e�e�e�g�l�G��H����J�N��W��e�e�e�d�g�m�G��I����W��^�D��w�u�u�u�u�l�G��I����W��^�D��e�e�d�e�f�m�U���Y���W��^�D��e�d�d�d�f�m�G��I����W��NךU���e�e�d�e�g�m�G��I����W��^�E��d�d�y�_�w�}�G��H����V��_�D��d�e�d�d�f�m�G��U���F�^�D��e�e�e�e�g�l�F��H����V��^��U���u�w�d�e�f�m�F��I����W��^�E��d�d�e�w�w�}�W���H����V��^�D��e�d�d�e�g�l�F��H���9F�L�E��e�e�d�d�g�l�F��H����V��_�D���_�u�u�e�g�m�G��H����V��^�E��e�e�d�d�f�q�}���Y����V��_�D��e�e�d�e�g�l�G��H����J�N��W��e�e�d�e�g�m�G��H����W��^�E��w�u�u�u�u�l�G��I����W��^�E��e�d�d�d�f�m�U���Y���W��^�E��d�d�d�e�f�l�G��H����V��NךU���e�e�e�e�g�l�F��I����W��_�D��e�d�y�_�w�}�G��H����V��_�E��d�e�d�d�g�l�G��U���F�_�D��e�d�d�e�f�m�F��H����W��_��U���u�w�e�d�f�l�F��I����V��^�D��e�e�e�w�w�}�W���I����V��_�D��e�e�d�e�f�m�F��I���9F�L�D��d�d�d�d�g�l�F��H����W��^�E���_�u�u�e�f�l�F��H����V��^�E��d�e�e�d�f�q�}���Y����W��_�D��d�e�d�d�g�l�F��I����J�N��W��d�e�e�d�f�l�F��I����W��_�E��w�u�u�u�u�m�F��H����W��^�D��e�d�d�d�f�l�U���Y���V��_�D��d�d�e�d�f�l�F��I����W��NךU���e�d�e�e�f�l�G��I����V��^�E��d�e�y�_�w�}�G��I����W��_�D��d�e�e�e�f�m�F��U���F�_�E��d�e�e�e�g�l�F��I����W��_��U���u�w�e�d�g�m�F��I����V��^�E��d�d�e�w�w�}�W���I����W��^�D��e�e�d�d�g�m�F��H���9F�L�D��e�d�d�e�g�m�F��H����W��^�E���_�u�u�e�f�l�F��I����V��_�E��e�e�d�d�f�q�}���Y����W��_�E��d�d�e�e�g�m�G��I����J�N��W��e�d�d�d�f�m�G��I����V��^�D��w�u�u�u�u�m�G��I����W��^�E��d�e�d�e�g�l�U���Y���V��^�E��d�e�e�d�g�l�F��H����V��NךU���e�d�d�d�g�l�G��I����W��^�D��e�d�y�_�w�}�G��H����V��^�E��e�e�e�e�f�m�G��U���F�_�D��d�e�e�e�f�m�F��I����V��^��U���u�w�e�e�f�m�F��I����W��^�E��d�e�e�w�w�}�W���I����W��^�E��e�e�d�d�g�l�F��I���9F�L�D��e�d�e�d�g�m�F��H����W��^�D���_�u�u�e�f�m�F��H����V��_�E��e�d�d�e�f�q�}���Y����V��^�E��e�d�d�d�g�m�G��H����J�N��W��e�e�d�e�g�l�F��I����V��_�D��w�u�u�u�u�m�G��I����V��_�E��d�e�d�d�g�l�U���Y���V��_�D��e�d�e�d�f�l�F��H����V��NךU���e�e�d�e�f�m�G��H����V��^�D��d�d�y�_�w�}�G��H����W��_�D��e�e�e�e�f�m�G��U���F�^�E��e�d�e�e�f�l�F��I����V��_��U���u�w�e�d�g�m�F��H����W��^�E��e�d�d�w�w�}�W���I����W��^�E��d�e�e�d�g�l�G��H���9F�L�E��e�e�e�d�g�m�F��I����W��_�E���_�u�u�e�g�m�F��H����W��^�E��e�e�d�d�g�q�}���Y����V��^�D��e�e�d�e�g�m�G��H����J�N��W��d�d�d�e�g�m�G��H����V��^�E��w�u�u�u�u�m�F��H����V��^�E��d�e�d�e�g�l�U���Y���V��^�D��e�d�d�d�f�m�F��H����W��NךU���e�e�e�e�f�m�F��I����V��^�D��e�e�y�_�w�}�G��I����V��^�D��d�e�e�e�f�m�G��U���F�^�D��d�e�e�d�g�l�G��I����V��_��U���u�w�e�e�f�m�G��H����W��^�E��d�d�e�w�w�}�W���I����W��_�E��d�e�e�d�g�m�F��I���9F�L�E��e�d�d�e�f�m�F��H����V��_�E���_�u�u�e�g�l�F��H����W��^�E��d�d�d�d�g�q�}���Y����W��_�D��d�d�d�d�g�l�F��H����J�N��W��e�e�d�d�g�m�F��I����W��_�E��w�u�u�u�u�m�G��I����W��^�E��e�d�d�d�f�m�U���Y���V��_�D��d�d�d�e�f�m�G��H����V��NךU���e�e�e�d�f�l�F��H����W��_�D��d�d�y�_�w�}�G��I����V��^�D��e�e�d�d�f�l�G��U���F�^�D��e�d�e�e�f�l�F��H����W��_��U���u�w�e�e�f�m�G��H����V��^�D��e�d�e�w�w�}�W���I����W��_�D��d�e�d�e�f�l�F��H���9F�L�E��d�e�d�d�f�m�G��I����W��_�D���_�u�u�e�g�m�G��H����V��^�E��e�e�d�d�f�q�}���Y����V��_�E��d�e�e�d�g�l�G��H����J�N��W��e�e�e�e�g�m�G��I����W��_�D��w�u�u�u�u�l�F��H����W��_�E��e�d�e�e�f�l�U���Y���W��_�E��d�e�d�e�f�m�G��I����W��NךU���d�d�d�e�f�l�F��I����V��_�E��d�e�y�_�w�}�F��H����W��^�D��e�e�d�d�f�l�G��U���F�_�D��e�d�e�d�f�l�F��H����V��_��U���u�w�d�d�g�l�F��H����W��^�E��d�e�d�w�w�}�W���H����V��^�D��e�e�d�e�g�l�G��I���9F�L�D��d�e�d�e�f�l�F��H����V��_�D���_�u�u�d�f�l�G��H����V��^�E��d�e�d�d�f�q�}���Y����W��_�D��d�d�e�e�g�l�F��I����J�N��W��d�e�e�e�f�l�G��H����W��_�E��w�u�u�u�u�l�F��H����W��_�D��e�e�d�e�g�m�U���Y���W��_�E��e�d�e�e�f�l�G��H����V��NךU���d�d�e�d�f�m�G��I����V��^�D��e�d�y�_�w�}�F��I����W��^�E��d�e�d�e�f�m�G��U���F�_�D��d�d�e�e�g�l�G��H����V��^��U���u�w�d�d�f�m�F��I����W��^�D��d�d�e�w�w�}�W���H����V��_�D��d�e�e�e�f�l�G��H���9F�L�D��e�e�e�d�f�m�G��H����W��^�D���_�u�u�d�f�m�F��I����W��_�E��d�d�d�d�g�q�}���Y����V��^�E��d�d�d�e�g�m�F��H����J�N��W��d�e�e�d�g�m�G��I����V��^�D��w�u�u�u�u�l�F��I����V��_�D��e�d�e�e�g�l�U���Y���W��^�E��d�d�d�d�f�m�G��H����W��NךU���d�d�e�e�f�l�F��I����W��_�E��e�e�y�_�w�}�F��I����W��_�D��e�e�e�e�g�m�G��U���F�_�E��e�d�e�d�g�m�F��I����V��_��U���u�w�d�d�g�m�F��H����W��^�D��d�d�e�w�w�}�W���H����V��_�D��e�e�d�e�f�m�G��I���9F�L�D��e�e�e�e�g�m�G��I����W��_�E���_�u�u�d�f�m�G��I����V��^�E��d�d�e�e�g�q�}���Y����W��_�E��d�d�e�d�g�m�F��H����J�N��W��e�d�d�e�f�m�F��H����V��_�E��w�u�u�u�u�l�G��H����V��_�D��e�e�e�e�f�l�U���Y���W��_�E��d�e�d�e�f�l�G��I����V��NךU���d�d�d�d�g�m�F��I����W��^�D��d�e�y�_�w�}�F��H����W��_�E��d�e�e�e�f�l�G��U���F�_�D��e�d�d�e�f�l�G��I����W��^��U���u�w�d�e�f�l�G��I����W��^�E��e�d�e�w�w�}�W���H����V��_�D��e�d�e�e�g�m�F��I���9F�L�D��d�d�d�e�g�l�G��I����V��^�E���_�u�u�d�f�l�F��H����V��^�E��e�e�e�e�f�q�}���Y����W��_�D��d�e�d�d�f�l�F��H����J�N��W��e�d�e�d�f�l�G��H����W��_�D��w�u�u�u�u�l�G��I����W��^�D��d�d�d�d�f�m�U���Y���W��_�E��d�e�e�e�f�m�F��H����W��NךU���d�d�d�d�g�m�F��I����W��_�D��d�d�y�_�w�}�F��H����W��_�E��e�d�d�d�f�l�F��U���F�_�D��d�e�e�d�f�l�F��H����W��_��U���u�w�d�e�f�l�F��I����V��_�D��e�d�e�w�w�}�W���H����W��^�E��e�e�d�d�f�l�F��I���9F�L�D��d�d�d�d�f�m�G��I����W��_�E���_�u�u�d�f�l�F��I����V��_�D��e�e�d�d�f�q�}���Y����V��^�E��e�e�d�d�f�l�G��I����J�N��W��d�e�e�e�f�m�F��H����W��^�E��w�u�u�u�u�l�F��I����V��_�E��d�d�e�d�f�m�U���Y���W��^�D��d�e�d�d�g�l�F��I����W��NךU���d�d�e�e�f�m�G��H����V��_�E��e�d�y�_�w�}�F��I����V��_�E��d�d�d�e�g�m�G��U���F�_�E��d�e�d�d�g�m�F��H����V��^��U���u�w�d�d�g�l�G��H����V��_�E��d�e�e�w�w�}�W���H����W��_�E��e�e�e�d�g�l�G��H���9F�L�D��d�e�e�d�f�m�G��I����W��^�E���_�u�u�d�f�m�F��H����V��^�D��d�e�d�e�f�q�}���Y����V��_�D��d�d�d�e�f�l�F��H����J�N��W��d�e�d�e�g�m�G��I����W��^�D��w�u�u�u�u�l�F��H����V��^�E��d�e�e�d�f�m�U���Y���W��^�D��e�e�e�d�f�m�F��I����W��NךU���d�d�e�d�f�l�F��I����V��^�D��d�d�y�_�w�}�F��I����V��^�D��e�d�d�d�f�m�F��U���F�_�D��e�e�e�d�f�m�G��H����W��_��U���u�w�d�d�f�l�G��I����W��_�E��d�d�d�w�w�}�W���H����W��^�E��e�d�e�d�g�m�G��H���9F�L�D��e�d�d�d�g�l�G��I����V��^�E���_�u�u�d�f�m�F��I����V��^�D��d�e�e�d�f�q�}���Y����V��^�D��d�d�d�e�f�l�G��H����J�N��W��d�d�e�d�f�l�F��H����W��_�E��w�u�u�u�u�l�F��H����V��_�E��d�e�d�d�f�l�U���Y���W��_�D��e�e�d�e�f�m�F��H����W��NךU���d�d�d�e�g�m�F��I����W��^�D��e�d�y�_�w�}�F��H����W��_�D��d�d�d�e�f�l�F��U���F�_�E��d�d�d�d�f�m�F��H����W��^��U���u�w�d�d�g�l�G��I����W��_�E��e�d�e�w�w�}�W���H����W��^�D��d�d�d�d�g�l�G��I���9F�L�D��d�e�e�d�f�m�G��I����W��^�D���_�u�u�d�f�l�F��H����W��_�D��e�d�e�e�f�q�}���Y����W��_�D��d�e�e�d�f�l�G��I����J�N��W��d�e�d�d�g�m�F��H����W��_�E��w�u�u�u�u�l�F��H����V��^�E��d�e�d�e�g�l�U���Y���W��_�E��e�e�d�e�f�m�F��H����W��NךU���d�d�d�e�g�l�F��I����V��^�D��d�d�y�_�w�}�F��H����V��_�E��d�d�d�e�f�m�G��U���F�_�D��d�e�d�d�g�l�G��H����V��_��U���u�w�d�d�f�l�G��I����V��_�E��e�e�e�w�w�}�W���H����V��_�E��d�e�e�d�g�l�G��I���9F�L�D��d�e�d�e�g�l�F��I����W��_�E���_�u�u�d�f�l�F��I����W��^�D��e�d�e�e�f�q�}���Y����W��^�D��e�d�e�e�f�l�G��I����J�N��W��d�d�d�e�f�l�G��H����W��_�D��w�u�u�u�u�m�G��I����V��^�E��d�e�d�d�f�m�U���Y���V��^�E��d�d�d�d�f�l�F��I����V��NךU���e�e�e�e�f�l�F��H����W��^�E��e�e�y�_�w�}�G��I����V��^�E��d�d�d�d�g�l�F��U���F�^�E��d�d�e�e�g�l�F��H����W��_��U���u�w�e�e�g�l�F��I����V��_�E��d�d�d�w�w�}�W���I����V��^�D��d�d�d�d�g�m�F��H���9F�L�E��d�d�e�e�f�m�F��H����V��^�D���_�u�u�e�g�m�F��I����V��^�D��d�d�d�e�g�q�}���Y����V��^�E��d�e�d�e�f�l�F��H����J�N��W��e�e�d�e�g�m�G��H����W��_�D��w�u�u�u�u�m�G��H����V��_�E��d�e�e�d�f�l�U���Y���V��_�E��d�d�d�d�f�l�F��H����W��NךU���e�e�e�e�g�l�F��H����W��^�E��e�d�y�_�w�}�G��I����W��_�D��d�d�d�d�g�m�G��U���F�^�D��e�e�e�e�f�l�G��H����W��_��U���u�w�e�e�f�l�F��H����W��_�E��e�d�d�w�w�}�W���I����W��^�D��e�e�d�d�g�l�G��H���9F�L�E��e�d�e�d�f�m�G��H����W��_�E���_�u�u�e�g�m�F��I����W��^�D��d�d�d�d�g�q�}���Y����V��^�E��e�e�e�e�f�l�G��H����J�N��W��e�d�e�e�g�m�G��I����W��^�E��w�u�u�u�u�m�G��I����V��_�D��d�d�e�d�g�m�U���Y���V��_�D��d�e�d�d�f�m�F��I����W��NךU���e�e�e�d�g�l�F��H����V��_�D��e�e�y�_�w�}�G��I����W��^�E��e�d�d�e�f�m�F��U���F�^�D��e�d�e�e�g�m�G��H����V��_��U���u�w�e�e�f�l�G��H����V��_�D��e�e�e�w�w�}�W���I����W��^�E��e�d�d�d�f�l�F��I���9F�L�E��e�e�e�e�g�m�G��I����W��_�D���_�u�u�e�g�l�G��H����V��^�D��e�d�e�d�f�q�}���Y����W��^�D��e�d�e�d�f�l�G��I����J�N��W��e�e�e�d�f�m�F��H����W��_�E��w�u�u�u�u�m�G��I����V��_�D��d�d�e�e�f�l�U���Y���V��^�D��e�d�e�d�f�l�F��I����V��NךU���e�e�d�e�f�m�G��I����V��_�E��d�e�y�_�w�}�G��H����W��_�E��d�d�d�d�f�m�G��U���F�^�E��d�d�e�d�g�l�F��H����W��^��U���u�w�e�e�g�l�G��H����V��_�D��d�e�e�w�w�}�W���I����W��_�E��d�d�e�d�f�l�G��I���9F�L�E��e�e�d�d�f�m�F��I����W��_�E���_�u�u�e�g�l�G��H����W��_�D��d�e�e�e�f�q�}���Y����W��^�D��e�d�e�d�f�l�F��H����J�N��W��e�e�d�d�g�m�G��H����W��_�E��w�u�u�u�u�m�G��H����W��_�E��d�d�d�d�g�l�U���Y���V��^�E��e�d�d�e�g�m�F��H����V��NךU���e�e�d�e�g�m�G��I����V��^�E��d�e�y�_�w�}�G��H����V��^�D��d�e�e�e�g�l�F��U���F�^�E��e�d�e�d�f�m�G��I����W��_��U���u�w�e�e�g�l�G��I����V��^�E��e�e�e�w�w�}�W���I����W��^�E��e�e�e�e�g�m�G��H���9F�L�E��e�e�e�d�f�m�F��I����V��_�E���_�u�u�e�g�l�G��I����V��^�E��e�d�d�e�f�q�}���Y����W��_�D��e�e�d�e�g�m�G��I����J�N��W��e�e�e�d�g�l�F��H����V��^�D��w�u�u�u�u�m�G��I����V��_�E��e�e�d�d�f�m�U���Y���V��^�D��d�d�e�e�g�m�G��H����V��NךU���e�e�d�e�f�l�G��H����W��^�D��d�e�y�_�w�}�G��H����V��^�D��e�e�e�e�f�l�F��U���F�^�E��d�e�d�d�f�l�F��I����V��_��U���u�w�e�e�g�m�F��I����V��^�E��d�d�d�w�w�}�W���I����V��^�D��e�e�e�e�g�m�G��I���9F�L�E��e�e�e�e�g�m�G��I����V��^�E���_�u�u�e�g�m�F��H����W��^�E��d�e�e�d�g�q�}���Y����V��_�D��e�d�e�d�g�m�F��H����J�N��W��e�d�d�e�f�m�G��I����V��^�D��w�u�u�u�u�m�G��H����V��_�E��e�e�e�e�f�l�U���Y���V��_�E��d�d�d�d�g�m�G��I����W��NךU���e�e�e�d�g�m�G��I����W��^�D��e�e�y�_�w�}�G��I����W��^�D��e�e�e�d�f�m�F��U���F�^�D��e�d�d�d�f�l�F��I����W��_��U���u�w�e�e�f�m�G��H����W��^�E��e�e�e�w�w�}�W���I����V��_�E��d�d�d�e�g�l�G��H���9F�L�E��d�e�d�e�f�m�G��H����W��^�E���_�u�u�e�g�m�G��H����V��^�E��d�e�d�d�f�q�}���Y����V��_�D��d�d�d�e�g�m�F��I����J�N��W��e�d�d�e�g�l�G��I����V��^�D��w�u�u�u�u�m�G��H����W��_�D��e�e�d�d�g�m�U���Y���V��_�E��e�d�d�e�g�m�G��H����W��NךU���e�e�e�e�f�m�F��H����W��^�D��e�e�y�_�w�}�G��I����W��^�D��d�e�e�d�f�m�F��U���F�^�D��d�e�d�e�f�l�G��I����V��_��U���u�w�e�e�f�m�G��I����W��^�E��e�e�e�w�w�}�W���I����W��_�D��e�e�e�e�g�l�G��I���9F�L�E��d�d�d�d�g�l�G��H����W��_�E���_�u�u�e�g�m�F��I����V��_�E��d�d�d�e�f�q�}���Y����V��^�E��d�e�d�d�g�m�F��H����J�N��W��e�e�d�e�g�m�F��I����V��_�E��w�u�u�u�u�m�G��I����W��^�D��e�e�d�d�g�l�U���Y���V��^�D��e�e�e�d�f�m�G��H����W��NךU���e�e�e�d�g�m�G��H����V��^�D��d�e�y�_�w�}�G��I����V��^�E��e�e�e�d�f�m�F��U���F�^�E��d�d�e�d�f�m�F��I����V��^��U���u�w�e�e�g�l�G��H����V��^�E��d�e�d�w�w�}�W���I����W��^�D��d�d�e�e�g�l�F��H���9F�L�E��e�e�d�e�f�m�F��H����W��^�E���_�u�u�e�g�m�G��H����V��_�E��d�d�d�d�g�q�}���Y����V��_�E��d�d�e�e�g�m�F��H����J�N��W��e�e�e�d�f�l�G��H����V��_�D��w�u�u�u�u�m�G��I����V��^�D��e�e�d�e�g�m�U���Y���V��^�E��e�e�e�e�g�m�G��H����V��NךU���d�d�d�d�f�m�G��I����V��^�D��d�d�y�_�w�}�F��H����V��^�D��d�e�e�d�f�m�G��U���F�_�D��d�d�d�e�f�m�G��I����V��_��U���u�w�d�d�f�l�G��H����V��^�E��d�d�d�w�w�}�W���H����V��^�D��d�e�e�e�g�l�F��I���9F�L�D��d�d�d�d�f�l�F��H����W��^�E���_�u�u�d�f�l�F��H����W��^�E��d�e�e�e�f�q�}���Y����W��^�E��e�e�e�e�g�m�F��I����J�N��W��d�d�e�e�f�m�G��I����V��^�D��w�u�u�u�u�l�F��H����W��_�E��e�e�d�e�g�m�U���Y���W��_�D��d�d�e�e�f�l�G��H����V��NךU���d�d�d�e�g�l�F��I����W��^�E��d�d�y�_�w�}�F��H����V��^�D��e�e�e�d�f�l�F��U���F�_�D��e�d�d�d�g�m�F��I����W��_��U���u�w�d�d�f�m�F��I����V��^�E��d�d�d�w�w�}�W���H����V��^�D��d�d�e�e�g�m�F��I���9F�L�D��e�d�e�d�f�m�G��I����V��^�D���_�u�u�d�f�l�G��H����W��^�E��d�d�e�d�f�q�}���Y����W��^�E��d�d�e�d�g�m�F��I����J�N��W��d�d�e�e�g�m�G��I����V��^�D��w�u�u�u�u�l�F��H����W��^�D��e�e�e�d�f�m�U���Y���W��^�D��d�e�e�d�g�m�G��I����W��NךU���d�d�d�d�f�l�G��I����V��^�E��e�e�y�_�w�}�F��H����V��_�D��e�e�e�d�g�m�F��U���F�_�E��d�d�e�d�f�l�G��I����V��_��U���u�w�d�d�g�l�F��H����V��^�E��d�e�e�w�w�}�W���H����W��_�D��d�e�d�e�g�l�F��H���9F�L�D��d�e�e�d�g�m�F��H����W��_�E���_�u�u�d�f�l�F��I����V��^�E��e�d�d�e�g�q�}���Y����W��_�E��d�d�e�e�g�m�G��I����J�N��W��d�e�e�d�f�m�G��H����V��^�D��w�u�u�u�u�l�F��I����W��_�D��e�e�d�d�f�m�U���Y���W��^�D��d�e�e�e�g�l�G��H����V��NךU���d�d�d�d�f�m�G��H����W��^�E��d�d�y�_�w�}�F��H����V��^�E��d�e�e�e�g�m�G��U���F�_�E��d�d�d�d�g�l�G��I����W��^��U���u�w�d�d�g�m�F��H����V��^�E��d�e�e�w�w�}�W���H����V��_�D��e�e�e�e�g�m�F��H���9F�L�D��d�e�e�d�f�l�F��H����V��^�D���_�u�u�d�f�l�F��I����W��_�E��e�d�e�e�g�q�}���Y����W��^�D��e�d�d�d�g�m�G��H����J�N��W��d�e�e�e�f�m�G��H����V��^�E��w�u�u�u�u�l�F��I����V��_�D��e�e�e�d�g�l�U���Y���W��^�E��e�e�d�e�g�m�G��I����V��NךU���d�d�d�d�g�l�F��I����W��^�E��d�d�y�_�w�}�F��H����W��_�D��d�e�e�e�g�m�G��U���F�_�E��e�d�e�e�f�m�G��H����W��_��U���u�w�d�d�g�m�G��I����V��_�D��d�d�d�w�w�}�W���H����V��_�D��e�e�e�d�f�l�G��H���9F�L�D��d�e�d�d�g�m�G��H����W��^�E���_�u�u�d�f�l�F��I����V��^�D��d�d�e�d�f�q�}���Y����W��^�E��e�e�e�d�f�l�F��H����J�N��W��d�e�e�d�f�l�G��I����W��^�E��w�u�u�u�u�l�F��I����V��_�E��d�d�d�d�g�l�U���Y���W��^�E��d�d�e�d�f�m�F��H����W��NךU���d�d�d�d�g�l�F��I����V��_�E��e�d�y�_�w�}�F��H����V��_�E��d�d�d�d�g�m�F��U���F�_�E��e�d�d�e�g�m�F��H����W��^��U���u�w�d�d�g�m�G��H����W��_�D��d�e�d�w�w�}�W���H����V��^�E��d�e�d�d�f�m�F��I���9F�L�D��d�d�e�e�g�l�F��H����V��_�D���_�u�u�d�f�l�F��H����W��^�D��d�d�d�d�g�q�}���Y����W��^�E��e�d�d�e�f�l�F��I����J�N��W��d�e�d�e�f�l�F��I����W��_�E��w�u�u�u�u�l�F��H����V��_�E��d�d�e�d�f�m�U���Y���W��^�E��d�e�d�e�g�m�F��I����V��NךU���d�d�d�d�g�l�G��I����V��_�E��d�e�y�_�w�}�F��H����W��_�E��e�d�d�d�g�m�F��U���F�_�E��e�d�d�e�g�l�F��H����W��_��U���u�w�d�d�g�l�G��I����W��_�D��e�e�d�w�w�}�W���H����W��_�D��d�d�e�d�f�m�G��H���9F�L�D��d�d�d�e�f�m�G��H����V��_�D���_�u�u�d�f�l�G��I����W��_�D��d�e�e�e�f�q�}���Y����W��^�D��e�d�e�e�f�l�G��H����J�N��W��d�d�e�d�f�l�F��H����W��_�E��w�u�u�u�u�l�F��I����V��^�E��d�d�d�d�g�l�U���Y���W��_�D��d�d�d�e�g�m�F��H����V��NךU���d�d�d�e�f�l�F��I����W��_�D��e�d�y�_�w�}�F��H����W��^�D��d�d�d�e�f�m�F��U���F�_�D��e�e�d�d�f�m�F��H����V��^��U���u�w�d�d�f�l�G��I����W��_�D��e�d�e�w�w�}�W���H����W��^�D��d�d�d�d�f�l�G��I���9F�L�D��e�e�d�e�g�m�F��H����W��^�E���_�u�u�d�f�l�G��I����W��_�D��e�d�d�d�g�q�}���Y����W��_�D��d�d�e�d�f�l�G��H����J�N��W��d�d�d�d�g�l�F��H����W��_�D��w�u�u�u�u�l�F��I����W��^�D��d�d�d�e�f�l�U���Y���W��_�E��e�d�d�d�f�m�F��H����V��NךU���d�d�d�d�g�m�F��I����W��_�D��e�d�y�_�w�}�F��H����V��^�E��e�d�d�e�f�m�G��U���F�_�D��e�e�d�e�f�m�G��H����V��^��U���u�w�d�d�f�m�F��H����W��_�D��e�d�d�w�w�}�W���H����V��_�E��e�d�d�d�f�l�G��H���9F�L�D��d�e�e�d�f�m�G��I����W��_�E���_�u�u�d�f�l�F��I����W��_�D��e�d�e�e�f�q�}���Y����W��^�E��e�e�e�e�f�l�G��I����J�N��W��d�d�d�e�g�l�G��H����W��_�D��w�u�u�u�u�l�F��H����W��^�E��d�d�d�e�f�l�U���Y���W��_�D��d�d�e�d�f�m�F��H����V��NךU���e�e�e�e�g�m�G��I����V��_�D��e�d�y�_�w�}�G��I����W��^�D��e�d�d�e�f�l�F��U���F�^�E��d�e�e�e�g�m�G��H����W��_��U���u�w�e�e�g�m�F��H����W��_�D��e�d�e�w�w�}�W���I����V��_�D��e�d�e�d�f�l�G��H���9F�L�E��e�d�d�e�f�m�F��H����W��^�D���_�u�u�e�g�m�G��I����W��^�D��e�d�e�d�f�q�}���Y����V��_�D��e�d�e�d�f�l�G��I����J�N��W��e�e�d�e�f�l�G��I����W��_�D��w�u�u�u�u�m�G��H����W��_�D��d�d�d�d�g�m�U���Y���V��^�E��e�e�d�d�f�m�F��H����V��NךU���e�e�e�e�f�m�G��I����W��_�D��d�d�y�_�w�}�G��I����W��^�D��e�d�d�d�g�m�G��U���F�^�E��e�d�d�d�f�m�F��H����V��^��U���u�w�e�e�g�l�F��H����V��_�D��e�d�d�w�w�}�W���I����W��_�D��d�e�d�d�f�m�G��I���9F�L�E��d�e�e�d�g�l�G��H����V��_�E���_�u�u�e�g�m�F��H����W��^�D��d�e�e�e�g�q�}���Y����V��^�E��d�e�d�d�f�l�F��I����J�N��W��e�e�e�d�g�m�G��I����W��^�D��w�u�u�u�u�m�G��I����V��^�E��d�d�e�d�g�m�U���Y���V��^�D��d�e�e�d�g�l�F��I����W��NךU���e�e�e�d�f�l�G��I����W��_�D��e�d�y�_�w�}�G��I����V��_�E��d�d�d�d�f�m�G��U���F�^�E��d�e�e�d�g�l�F��H����W��^��U���u�w�e�e�g�m�F��H����W��_�D��e�e�d�w�w�}�W���I����W��^�D��d�d�d�d�f�m�G��H���9F�L�E��d�e�e�d�g�l�F��H����V��^�E���_�u�u�e�g�m�F��H����V��^�D��d�d�e�d�g�q�}���Y����V��^�E��d�d�e�d�f�l�F��H����J�N��W��e�e�d�d�f�m�F��I����W��_�D��w�u�u�u�u�m�G��H����V��_�D��d�d�d�e�g�m�U���Y���V��^�E��d�d�e�e�g�m�F��H����V��NךU���e�e�e�d�g�l�F��H����W��_�E��d�d�y�_�w�}�G��I����V��^�E��e�d�d�d�g�l�F��U���F�^�E��e�d�d�e�f�m�G��H����V��_��U���u�w�e�e�g�l�G��H����W��_�D��d�d�e�w�w�}�W���I����W��^�E��e�e�d�d�f�l�F��I���9F�L�E��d�d�d�e�g�m�G��I����W��_�E���_�u�u�e�g�m�F��H����W��^�D��d�d�e�d�g�q�}���Y����V��_�D��d�d�e�d�f�l�F��I����J�N��W��e�e�d�d�g�m�F��I����W��_�E��w�u�u�u�u�m�G��H����W��_�E��d�d�d�e�f�l�U���Y���V��^�D��d�d�d�d�g�l�F��H����W��NךU���e�e�e�d�f�m�F��H����W��_�D��d�e�y�_�w�}�G��I����V��_�E��d�d�d�d�f�l�F��U���F�^�E��d�e�d�e�g�m�F��H����W��^��U���u�w�e�e�g�l�F��H����W��^�E��e�e�d�w�w�}�W���I����W��^�E��d�d�e�e�g�m�G��I���9F�L�E��d�d�e�d�g�l�G��H����V��^�D���_�u�u�e�g�m�F��I����W��_�E��e�e�d�d�f�q�}���Y����V��_�E��d�d�d�d�g�m�G��I����J�N��W��e�e�d�e�f�l�G��H����V��^�D��w�u�u�u�u�m�G��H����W��^�D��e�e�e�d�g�l�U���Y���V��^�D��d�d�d�e�g�m�G��I����W��NךU���e�e�e�d�f�l�G��I����W��^�D��e�d�y�_�w�}�G��I����V��^�D��e�e�e�e�f�m�G��U���F�^�E��e�d�e�d�g�l�G��I����V��_��U���u�w�e�e�g�l�G��I����V��^�E��e�e�e�w�w�}�W���I����W��_�E��d�d�e�e�g�m�G��I���9F�L�E��d�e�d�e�g�m�F��I����V��^�E���_�u�u�e�g�m�F��H����V��^�E��e�d�e�e�g�q�}���Y����V��^�D��e�d�e�e�g�m�G��I����J�N��W��e�e�d�d�g�l�F��H����V��_�E��w�u�u�u�u�m�G��H����V��_�D��e�e�e�d�f�l�U���Y���V��^�E��d�e�e�d�g�l�G��H����V��NךU���e�e�e�d�g�m�G��H����V��^�E��d�d�y�_�w�}�G��I����V��_�D��d�e�e�e�g�m�G��U���F�^�E��d�d�d�e�g�m�F��I����V��_��U���u�w�e�e�g�m�F��I����V��^�E��e�e�e�w�w�}�W���I����V��^�D��d�e�d�e�g�l�G��I���9F�L�E��d�d�d�d�f�m�F��H����W��_�E���_�u�u�e�g�m�F��H����W��_�E��e�e�e�e�g�q�}���Y����V��_�D��e�e�d�d�g�m�G��I����J�N��W��e�e�e�d�f�l�F��I����V��^�D��w�u�u�u�u�m�G��I����W��_�E��e�e�d�d�f�m�U���Y���V��^�E��e�e�e�d�f�m�G��H����V��NךU���e�e�e�d�g�l�F��H����W��^�E��d�e�y�_�w�}�G��I����W��_�D��e�e�e�e�g�l�F��U���F�^�E��e�e�d�e�g�m�F��I����W��^��U���u�w�e�e�g�l�F��H����V��^�E��d�d�e�w�w�}�W���I����W��_�E��e�e�e�e�g�l�F��H���9F�L�E��e�d�e�e�g�l�G��H����W��^�D���_�u�u�e�g�m�G��H����V��^�E��e�d�e�e�f�q�}���Y����V��_�D��d�e�d�d�g�m�G��I����J�N��W��e�e�d�d�f�m�G��I����V��_�E��w�u�u�u�u�m�G��H����V��_�D��e�e�d�e�f�m�U���Y���V��^�E��d�e�d�d�g�m�G��H����V��NךU���e�e�e�e�g�l�F��I����V��^�D��e�e�y�_�w�}�G��I����V��_�E��e�e�e�e�f�m�G��U���F�^�E��d�d�d�e�g�m�F��I����V��^��U���u�w�e�e�g�m�F��I����W��^�E��e�d�e�w�w�}�W���I����V��^�E��e�d�d�e�g�l�G��I���9F�L�E��e�d�d�e�g�m�G��H����W��_�E���_�u�u�e�g�m�G��I����W��_�E��e�d�e�d�g�q�}���Y����V��^�D��d�e�d�d�g�m�G��I����J�N��W��e�e�e�d�g�m�F��I����V��_�D��w�u�u�u�u�m�G��I����V��^�E��e�e�d�e�f�l�U���Y���V��^�E��e�e�d�d�g�m�G��H����V��NךU���e�e�e�e�g�m�F��H����V��^�D��d�d�y�_�w�}�G��I����V��^�E��e�e�e�e�f�m�F��U���F�_�D��d�e�d�d�f�l�F��I����V��^��U���u�w�d�d�f�l�F��H����W��^�E��e�e�d�w�w�}�W���H����W��_�D��d�d�e�e�g�l�G��I���9F�L�D��d�d�e�d�f�m�F��I����W��_�E���_�u�u�d�f�l�F��I����W��^�E��e�e�d�d�g�q�}���Y����W��^�D��e�d�e�d�g�m�G��H����J�N��W��d�d�d�d�f�m�F��H����V��^�E��w�u�u�u�u�l�F��H����V��^�D��e�e�d�d�g�m�U���Y���W��_�E��d�e�e�d�g�l�G��H����V��NךU���d�d�d�d�g�m�G��H����V��^�E��d�d�y�_�w�}�F��H����V��_�E��d�e�e�e�g�m�G��U���F�_�D��d�e�d�d�g�l�G��I����V��_��U���u�w�d�d�f�m�F��I����V��^�E��d�e�d�w�w�}�W���H����V��^�E��d�e�d�e�g�l�G��H���9F�L�D��d�d�d�e�g�l�F��H����W��_�D���_�u�u�d�f�l�F��I����V��^�E��e�e�d�e�g�q�}���Y����W��_�E��e�e�d�d�g�m�G��H����J�N��W��d�d�e�d�f�m�G��H����V��^�D��w�u�u�u�u�l�F��I����V��_�E��e�e�d�e�f�l�U���Y���W��_�E��d�e�d�e�g�l�G��H����W��NךU���d�d�d�d�g�m�F��I����W��^�E��e�e�y�_�w�}�F��H����W��^�E��e�e�e�e�f�l�F��s���K�\-�����8�'�d�_�w�}�L���Y���P	��C��U���"�&��0�1�3��������~'��T�����0�u�h�_�w�}�Zӵ�����p	��Q'�����'�=�&��e�W�W���@��ƹF�R��9���&��0�3�9�8�1�������pT�N��N���6�;�!�;�w���������U/��R�����&��g�o�>�)����C��ƹF�R�����&��0�3�9�8�1�������pT�N��G��_�u�u�x�x���������U/��R�����&��g�_�w�}�}�������]��t�����:�,�u�u���A���C���F�C��6���3�0�:�,�i�}�W�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��d�e�d�d�f�l�F��H���F�^�E��e�e�e�e�g�l�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�d�d�g�m�G��I����V�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��^�E��d�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�F��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��d�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�l�F��I����V��^�W���u�u�w�e�g�m�G��I����W��_�E��e�e�e�e�u�}�W���[����V��^�E��e�e�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�d�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�D��d�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�f�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�d�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�f�m�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�l�F��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�e�u�}�W���[����W��_�D��d�e�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��H����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�g�l�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��d�d�e�e�g�m�G��I���F�_�D��d�d�d�d�f�l�G��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�e�u�}�W���[����W��_�D��e�e�e�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��I����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�e�e�f�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�g�m�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�E��e�d�e�e�g�m�G��I���F�_�D��d�d�d�d�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�e�u�}�W���[����W��_�D��d�e�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��H����V��^�E��y�_�u�u�f�l�F��H����W��_�D��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�e�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�f�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�E��d�d�e�e�g�m�G��I���F�_�D��d�d�d�d�g�l�F��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�e�u�}�W���[����W��_�D��e�d�d�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��H����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�e�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��^�E��d�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�f�l�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�d�d�d�f�l�F��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�e�u�}�W���[����W��_�D��d�e�d�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�e�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�f�m�F��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�D��d�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�F��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�D��d�e�e�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�e�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�g�l�F��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�D��d�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�d�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�f�l�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�E��d�e�e�e�g�m�G��I���F�_�D��d�d�d�d�g�m�G��H����W��_�W���u�u�w�d�f�l�F��H����V��^�D��d�d�d�d�u�}�W���[����W��_�D��e�e�d�e�f�l�F��H����FǻN��D��d�d�d�d�f�l�G��I����W��_�D��y�_�u�u�f�l�F��H����W��_�D��d�d�d�d�f�l�[�ԜY���W��_�D��d�e�e�e�g�l�F��H����W�d��U���d�d�d�d�f�l�F��I����W��_�D��d�w�u�u�w��F��H����W��^�D��d�d�d�d�f�l�F���Y���D��_�D��d�d�d�d�g�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�d�y�]�}�W��H����W��_�D��e�d�d�d�f�l�F��H���F�_�D��d�d�d�d�f�m�G��H����W��_�W���u�u�w�d�f�l�F��H����W��^�D��d�d�d�d�u�}�W���[����W��_�D��e�e�d�e�f�l�F��H����FǻN��D��d�d�d�d�f�l�G��H����W��_�D��y�_�u�u�f�l�F��H����W��^�D��d�d�d�d�f�l�[�ԜY���W��_�D��d�d�e�d�f�l�F��H����W�d��U���d�d�d�d�f�l�F��H����W��_�D��d�w�u�u�w��G��I����V��^�E��e�d�d�d�f�l�F���Y���D��^�E��e�e�e�e�f�m�G��H����W��L����u�e�e�e�g�m�G��I����W��_�D��d�d�d�y�]�}�W��I����V��^�E��e�d�d�d�f�l�F��H���F�^�E��e�e�e�e�g�m�F��H����W��_�W���u�u�w�e�g�m�G��I����V��^�D��d�d�d�d�u�}�W���[����V��^�E��d�d�e�e�f�l�F��H����FǻN��E��e�e�e�e�g�m�G��H����W��_�D��y�_�u�u�g�m�G��I����V��_�E��d�d�d�d�f�l�[�ԜY���V��^�E��e�d�d�d�g�l�F��H����W�d��U���e�e�e�e�g�m�G��I����W��_�D��d�w�u�u�w��G��I����V��_�D��d�d�d�d�f�l�F���Y���D��^�E��e�e�e�d�g�l�F��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�d�d�y�]�}�W��I����V��^�E��d�e�d�d�f�l�F��H���F�^�E��e�e�e�e�g�l�F��H����W��_�W���u�u�w�e�g�m�G��I����V��^�D��d�d�d�d�u�}�W���[����V��^�E��d�d�e�d�f�l�F��H����FǻN��E��e�e�e�e�g�l�F��I����W��_�D��y�_�u�u�g�m�G��I����W��^�E��d�d�d�d�f�l�[�ԜY���V��^�E��e�d�e�d�f�l�F��H����W�d��U���e�e�e�e�g�m�G��H����W��_�D��d�w�u�u�w��G��I����V��_�E��d�d�d�d�f�l�F���Y���D��^�E��e�e�d�d�g�l�G��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�d�d�y�]�}�W��I����V��^�E��e�e�d�d�f�l�F��H���F�^�E��e�e�e�d�g�l�F��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�d�u�}�W���[����V��^�E��d�d�d�d�f�l�F��H����FǻN��E��e�e�e�e�g�m�F��I����W��_�D��y�_�u�u�g�m�G��I����V��^�E��d�d�d�d�f�l�[�ԜY���V��^�E��d�d�e�e�f�l�F��H����W�d��U���e�e�e�e�g�m�F��H����W��_�D��d�w�u�u�w��G��I����V��_�E��e�d�d�d�f�l�F���Y���D��^�E��e�e�e�d�f�l�F��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�d�d�y�]�}�W��I����V��^�D��d�d�d�d�f�l�F��H���F�^�E��e�e�e�d�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�d�u�}�W���[����V��^�E��e�d�e�d�f�l�F��H����FǻN��E��e�e�e�e�g�l�F��I����W��_�D��y�_�u�u�g�m�G��I����W��_�E��d�d�d�d�f�l�[�ԜY���V��^�E��d�e�d�d�f�l�F��H����W�d��U���e�e�e�e�g�m�F��H����W��_�D��d�w�u�u�w��G��I����V��_�E��e�d�d�d�f�l�F���Y���D��^�E��e�e�d�e�f�l�F��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�d�d�y�]�}�W��I����V��^�D��d�e�d�d�f�l�F��H���F�^�E��e�e�e�d�f�m�G��H����W��_�W���u�u�w�e�g�m�G��I����V��^�D��d�d�d�d�u�}�W���[����V��^�E��d�d�d�e�f�l�F��H����FǻN��E��e�e�e�e�g�l�F��H����W��_�D��y�_�u�u�g�m�G��I����W��^�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�d�d�d�g�l�F��H����W�d��U���e�e�e�e�g�m�F��H����V��^�E��e�w�u�u�w��G��I����V��^�E��d�e�e�e�g�m�G���Y���D��^�E��e�d�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����W��^�E��e�e�e�y�]�}�W��I����V��_�E��e�d�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�D��e�d�d�e�g�m�G��I����FǻN��E��e�e�e�e�f�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�d�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�d�d�f�m�G��I����V��L����u�e�e�e�g�m�G��H����W��^�E��e�e�d�y�]�}�W��I����V��^�D��e�e�e�e�g�m�G��H���F�^�E��e�e�e�d�f�m�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�d�d�d�g�m�G��I����FǻN��E��e�e�e�e�g�l�G��H����V��^�E��y�_�u�u�g�m�G��I����W��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�d�e�d�g�m�G��I����W�d��U���e�e�e�e�g�m�F��H����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�d�d�g�m�F��I����V��L����u�e�e�e�g�m�G��H����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�d�e�e�g�m�G��I���F�^�E��e�e�e�d�f�l�F��I����V��^�W���u�u�w�e�g�m�G��I����V��_�E��e�e�e�d�u�}�W���[����V��^�E��d�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�e�g�m�[�ԜY���V��^�E��d�e�d�e�g�m�G��I����V�d��U���e�e�e�e�g�m�F��H����V��^�E��d�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�F���Y���D��^�E��e�e�d�d�f�m�G��I����V��L����u�e�e�e�g�m�G��H����V��^�E��e�e�e�y�]�}�W��I����V��^�D��e�d�e�e�g�m�G��H���F�^�E��e�e�e�e�g�l�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�d�u�}�W���[����V��^�E��e�e�e�d�g�m�G��I����FǻN��E��e�e�e�e�g�m�F��H����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�l�[�ԜY���V��^�E��e�d�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�E��d�w�u�u�w��G��I����V��^�D��d�e�e�e�g�m�F���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�d�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�d�u�}�W���[����W��_�D��d�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��H����V��^�E��y�_�u�u�f�l�F��H����V��^�D��e�e�e�e�f�m�[�ԜY���W��_�D��d�e�e�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�f�m�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�d�e�y�]�}�W��H����W��_�E��e�e�e�e�g�m�G��I���F�_�D��d�d�d�e�f�l�F��I����V��_�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�e�u�}�W���[����W��_�D��d�e�d�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��I����V��^�D��y�_�u�u�f�l�F��H����W��_�D��e�e�e�e�f�m�[�ԜY���W��_�D��d�d�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�e�d�e�g�l�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�d�e�y�]�}�W��H����W��^�D��d�e�e�e�g�m�G��I���F�_�D��d�d�d�d�g�m�G��I����V��_�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�E��d�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�g�l�G��H����V��^�D��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�f�m�[�ԜY���W��_�D��e�e�d�e�g�m�G��I����W�d��U���d�d�d�d�f�l�G��H����V��^�E��d�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�F���Y���D��_�D��d�e�e�e�f�l�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�e�d�y�]�}�W��H����W��^�E��d�d�e�e�g�m�G��H���F�_�D��d�d�e�d�f�l�F��I����V��^�W���u�u�w�d�f�l�F��I����V��^�E��e�e�e�d�u�}�W���[����W��_�D��e�d�d�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��I����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�g�l�[�ԜY���W��_�D��d�e�e�d�f�m�G��I����W�d��U���d�d�d�d�f�m�F��H����V��^�E��d�w�u�u�w��F��H����V��_�D��d�e�e�e�g�m�F���Y���D��_�D��d�d�e�e�g�l�F��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�e�e�y�]�}�W��H����W��_�E��d�d�e�e�g�m�G��I���F�_�D��d�d�e�d�g�m�F��I����V��^�W���u�u�w�d�f�l�F��I����W��_�E��e�e�e�d�u�}�W���[����W��_�D��e�d�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��I����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�g�l�[�ԜY���W��_�D��e�d�e�d�f�m�G��I����W�d��U���d�d�d�d�f�m�G��I����V��^�E��e�w�u�u�w��F��H����V��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�f�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�d�e�e�f�l�G��I����V��^�W���u�u�w�d�f�l�F��I����W��^�E��e�e�e�e�u�}�W���[����W��_�D��e�e�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��H����V��^�E��y�_�u�u�f�l�F��H����W��_�E��d�d�d�d�f�l�[�ԜY���W��_�D��e�d�e�e�g�l�F��H����W�d��U���d�d�d�d�f�m�G��I����W��_�D��d�w�u�u�w��F��H����V��_�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�d�d�f�l�G��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�e�y�]�}�W��H����W��_�E��e�e�d�d�f�l�F��I���F�_�D��d�d�e�d�g�m�G��H����W��_�W���u�u�w�d�f�l�F��I����W��_�D��d�d�d�d�u�}�W���[����W��_�D��e�d�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�F��I����W��_�D��y�_�u�u�f�l�F��H����V��^�D��d�d�d�d�f�l�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����W�d��U���d�d�d�d�f�m�F��I����W��_�D��e�w�u�u�w��F��H����V��_�E��e�d�d�d�f�l�G���Y���D��_�D��d�d�d�e�f�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�e�y�]�}�W��H����W��^�E��e�d�d�d�f�l�F��I���F�_�D��d�d�d�e�g�l�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�e�u�}�W���[����W��_�E��e�e�d�e�f�l�F��H����FǻN��D��d�d�d�d�g�l�F��I����W��_�E��y�_�u�u�f�l�F��H����W��^�E��d�d�d�d�g�l�[�ԜY���W��_�D��e�d�d�e�f�l�F��H����W�d��U���d�d�d�d�f�l�F��I����W��_�D��d�w�u�u�w��F��H����W��_�D��e�d�d�d�f�l�F���Y���D��_�D��d�e�e�d�f�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�e�e�y�]�}�W��H����W��^�D��e�d�d�d�f�l�F��I���F�_�D��d�d�d�e�g�m�F��H����W��^�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�D��d�e�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�l�F��I����W��_�E��y�_�u�u�f�l�F��H����W��_�D��d�d�d�d�g�l�[�ԜY���W��_�D��d�e�d�d�g�l�F��H����W�d��U���d�d�d�d�f�l�F��I����W��_�D��e�w�u�u�w��F��H����W��^�D��e�d�d�d�f�l�G���Y���D��_�D��d�d�d�e�g�m�G��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�e�d�y�]�}�W��I����V��^�E��d�d�d�d�f�l�F��I���F�^�E��e�e�e�e�f�l�G��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�e�u�}�W���[����V��^�E��d�d�e�d�f�l�F��H����FǻN��E��e�e�e�e�g�m�F��I����W��_�E��y�_�u�u�g�m�G��I����V��_�D��d�d�d�d�g�m�[�ԜY���V��^�E��d�e�d�e�g�l�F��H����V�d��U���e�e�e�e�g�m�F��H����W��_�D��e�w�u�u�w��G��I����V��^�D��d�d�d�d�f�l�G���Y���D��^�E��e�d�d�e�g�m�G��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�e�e�y�]�}�W��I����V��_�E��d�d�d�d�f�l�F��I���F�^�E��e�e�e�d�f�m�G��H����W��^�W���u�u�w�e�g�m�G��I����V��_�D��d�d�d�e�u�}�W���[����V��^�D��e�e�d�d�f�l�F��H����FǻN��E��e�e�e�e�g�m�G��H����W��_�E��y�_�u�u�g�m�G��I����V��_�E��d�d�d�d�g�m�[�ԜY���V��^�E��e�e�d�d�f�l�F��H����V�d��U���e�e�e�e�g�l�G��I����W��_�D��e�w�u�u�w��G��I����W��^�E��d�d�d�d�f�l�G���Y���D��^�E��e�e�e�d�g�l�G��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�e�e�y�]�}�W��I����V��^�D��e�e�d�d�f�l�F��I���F�^�E��e�e�d�e�g�m�G��H����W��^�W���u�u�w�e�g�m�G��H����V��_�D��d�d�d�e�u�}�W���[����V��^�D��d�d�d�d�f�l�F��H����FǻN��E��e�e�e�e�f�l�F��I����W��_�E��y�_�u�u�g�m�G��I����V��^�E��d�d�d�d�g�m�[�ԜY���V��^�E��d�d�e�e�f�l�F��H����V�d��U���e�e�e�e�g�l�F��H����W��_�D��e�w�u�u�w��G��I����W��_�D��e�d�d�d�f�l�G���Y���D��^�E��d�e�e�e�g�l�G��H����W��L����u�e�e�e�g�m�F��I����W��_�D��d�e�d�y�]�}�W��I����V��^�E��e�e�d�d�f�l�F��H���F�^�E��e�e�e�e�g�l�F��H����W��^�W���u�u�w�e�g�m�G��I����V��^�D��d�d�d�d�u�}�W���[����V��^�E��e�d�d�e�f�l�F��H����FǻN��E��e�e�e�d�g�m�G��I����W��_�E��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�g�m�[�ԜY���V��^�E��d�e�e�e�f�l�F��H����V�d��U���e�e�e�e�g�m�F��I����W��_�D��d�w�u�u�w��G��I����V��_�E��e�d�d�d�f�l�F���Y���D��^�E��d�d�e�e�f�m�G��H����W��L����u�e�e�e�g�m�F��I����W��_�D��d�d�e�y�]�}�W��I����V��_�D��e�d�d�d�f�l�F��I���F�^�E��e�e�e�e�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�e�u�}�W���[����V��^�D��d�e�d�d�f�l�F��H����FǻN��E��e�e�e�d�f�l�G��H����W��_�D��y�_�u�u�g�m�G��I����W��^�D��d�d�d�d�f�l�[�ԜY���V��^�E��e�d�d�d�f�l�F��H����V�d��U���e�e�e�e�g�m�F��I����W��_�D��d�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�F���Y���D��^�E��d�d�e�e�f�l�G��H����W��L����u�e�e�e�g�m�F��I����W��_�D��d�d�d�y�]�}�W��I����V��_�E��e�d�d�d�f�l�F��H���F�^�E��e�e�e�d�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����V��_�E��e�e�e�e�u�}�W���[����V��^�D��d�e�d�e�g�m�G��I����FǻN��E��e�e�e�d�f�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�e�g�l�[�ԜY���V��^�E��d�e�e�d�f�m�G��I����V�d��U���e�e�e�e�g�m�G��H����V��^�E��d�w�u�u�w��G��I����V��_�E��d�e�e�e�g�m�F���Y���D��^�E��d�d�d�e�f�l�G��I����V��L����u�e�e�e�g�m�F��H����V��^�E��e�e�d�y�]�}�W��I����V��_�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�f�l�G��I����V��_�W���u�u�w�e�g�m�G��I����V��_�E��e�e�e�e�u�}�W���[����V��^�D��d�e�e�d�g�m�G��I����FǻN��E��e�e�e�d�g�l�F��H����V��^�D��y�_�u�u�g�m�G��I����W��_�E��e�e�e�e�f�m�[�ԜY���V��^�E��d�e�d�e�f�m�G��I����V�d��U���e�e�e�e�g�m�F��I����V��^�E��d�w�u�u�w��G��I����V��^�D��d�e�e�e�g�m�F���Y���D��^�E��d�e�d�d�g�l�G��I����V��L����u�e�e�e�g�m�F��H����V��^�E��e�e�e�y�]�}�W��I����V��^�D��e�d�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�F��I����V��^�W���u�u�w�e�g�m�G��H����V��^�E��e�e�d�e�u�}�W���[����V��^�D��e�d�d�d�g�m�G��H����FǻN��E��e�e�e�e�f�m�G��I����V��^�E��y�_�u�u�g�m�G��I����W��_�D��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�d�f�m�G��I����W�d��U���e�e�e�e�g�l�G��H����V��^�E��d�w�u�u�w��G��I����W��_�E��d�e�e�e�g�l�F���Y���D��^�E��e�e�d�e�f�m�F��I����W��L����u�e�e�e�g�m�G��I����V��^�E��e�d�e�y�]�}�W��I����V��^�D��d�e�e�e�g�m�G��I���F�^�E��e�e�d�e�f�l�G��I����V��_�W���u�u�w�e�g�m�G��H����V��^�E��e�e�d�e�u�}�W���[����V��^�D��d�e�e�e�g�m�G��H����FǻN��E��e�e�e�e�f�m�F��H����V��^�D��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�f�m�[�ԜY���V��^�E��e�d�d�e�f�m�G��I����V�d��U���e�e�e�e�g�m�F��I����V��^�E��d�w�u�u�w��G��I����V��_�D��e�e�e�e�g�l�F���Y���D��^�E��e�e�d�d�g�m�G��I����W��L����u�e�e�e�g�m�G��I����W��^�E��e�d�d�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�D��e�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��I����V��^�E��y�_�u�u�f�l�F��H����W��^�D��e�e�e�d�g�m�[�ԜY���W��_�D��d�e�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�G��H����V��^�E��e�w�u�u�w��F��H����V��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�g�l�F��I����V��L����u�d�d�d�f�l�F��H����V��^�E��d�e�d�y�]�}�W��H����W��_�D��d�e�e�e�g�m�F��H���F�_�D��d�d�e�d�f�m�G��I����V��^�W���u�u�w�d�f�l�F��I����W��_�E��e�e�e�e�u�}�W���[����W��_�E��e�e�d�d�g�m�G��I����FǻN��D��d�d�d�d�g�m�G��I����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�d�g�l�[�ԜY���W��_�D��d�d�e�e�g�m�G��I����W�d��U���d�d�d�d�f�l�G��H����V��^�E��e�w�u�u�w��F��H����W��^�E��d�e�e�e�g�m�G���Y���D��_�D��e�e�d�d�g�l�G��I����V��L����u�d�d�d�f�l�G��I����V��^�E��d�e�e�y�]�}�W��H����W��^�E��d�d�e�e�g�m�F��I���F�_�D��d�d�d�e�g�m�F��I����V��^�W���u�u�w�d�f�l�F��I����W��^�E��e�e�e�e�u�}�W���[����W��_�D��d�e�e�e�g�m�G��I����FǻN��D��d�d�d�e�f�l�F��I����V��^�D��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�f�l�[�ԜY���W��_�D��d�d�e�e�f�m�G��I����W�d��U���d�d�d�d�f�m�F��H����V��^�E��d�w�u�u�w��F��H����V��_�E��e�e�e�e�g�l�F���Y���D��_�D��e�e�e�d�g�l�F��I����W��L����u�d�d�d�f�l�G��I����V��^�E��e�d�e�y�]�}�W��H����W��_�E��e�d�e�e�g�m�G��H���F�_�D��d�e�d�d�g�l�F��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�e�d�e�u�}�W���[����W��^�D��d�e�e�e�g�m�G��H����FǻN��D��d�d�d�d�f�m�G��H����V��^�D��y�_�u�u�f�l�F��H����W��_�D��e�e�e�e�g�l�[�ԜY���W��_�E��d�d�e�e�f�m�G��I����W�d��U���d�d�d�d�g�l�F��H����V��^�E��d�w�u�u�w��F��H����W��_�E��e�e�e�e�g�l�F���Y���D��_�D��d�e�e�d�f�l�G��I����W��L����u�d�d�d�f�l�F��I����V��^�E��e�e�d�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�e�e�d�g�l�F��I����V��^�W���u�u�w�d�f�l�F��I����W��_�E��e�e�e�d�u�}�W���[����W��^�D��e�d�e�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��H����V��^�D��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�f�l�[�ԜY���W��_�E��e�d�d�e�g�m�G��I����W�d��U���d�d�d�d�g�m�G��H����V��^�E��e�w�u�u�w��F��H����V��^�E��d�e�e�e�g�m�F���Y���D��_�D��d�d�d�e�g�l�F��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�e�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��H���F�_�D��d�e�e�e�f�m�F��I����V��^�W���u�u�w�d�f�l�F��I����V��_�E��e�e�e�e�u�}�W���[����W��^�D��d�e�e�e�f�l�F��H����FǻN��D��d�d�d�d�f�m�F��H����W��_�D��y�_�u�u�f�l�F��H����W��^�E��d�d�d�d�f�m�[�ԜY���W��_�E��e�e�e�e�f�l�F��H����W�d��U���d�d�d�d�g�m�G��I����W��_�D��e�w�u�u�w��F��H����V��_�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�e�e�f�m�G��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�e�e�y�]�}�W��H����W��_�E��d�d�d�d�f�l�F��H���F�_�D��d�e�e�d�f�m�G��H����W��^�W���u�u�w�d�f�l�F��H����V��_�D��d�d�d�e�u�}�W���[����W��^�E��e�e�e�e�f�l�F��I����FǻN��D��d�d�d�d�g�l�F��I����W��_�D��y�_�u�u�f�l�F��H����W��^�D��d�d�d�d�f�l�[�ԜY���W��_�E��d�d�d�d�g�l�F��H����V�d��U���d�d�d�d�g�l�F��H����W��_�D��e�w�u�u�w��F��H����W��^�D��e�d�d�d�f�m�F���Y���D��_�D��d�d�d�e�f�m�F��H����V��L����u�d�d�d�f�l�F��I����W��_�D��d�e�d�y�]�}�W��H����W��_�D��d�e�d�d�f�l�F��H���F�_�D��d�e�d�d�f�l�F��H����W��^�W���u�u�w�d�f�l�F��I����V��^�D��d�d�d�d�u�}�W���[����W��_�E��e�d�d�d�f�l�F��H����FǻN��D��d�d�d�e�g�l�F��I����W��_�D��y�_�u�u�f�l�F��H����V��^�D��d�d�d�e�f�l�[�ԜY���W��_�D��e�d�d�e�f�l�F��H����V�d��U���d�d�d�d�f�m�F��H����W��_�D��e�w�u�u�w��F��H����W��^�D��e�d�d�d�f�l�F���Y���D��_�D��e�e�d�e�f�m�F��H����W��L����u�d�d�d�f�l�G��I����V��_�D��e�e�e�y�]�}�W��H����W��_�E��d�d�d�d�f�l�G��H���F�_�D��d�d�d�e�f�m�G��H����W��^�W���u�u�w�d�f�l�F��H����V��^�D��d�d�d�e�u�}�W���[����W��_�E��d�d�d�e�f�l�F��H����FǻN��D��d�d�d�d�g�m�F��H����W��_�D��y�_�u�u�f�l�F��H����V��^�D��d�d�d�e�f�m�[�ԜY���W��_�D��e�d�d�e�f�l�F��H����V�d��U���d�d�d�d�f�m�F��I����W��_�D��e�w�u�u�w��F��H����W��_�D��d�d�d�d�f�m�G���Y���D��_�D��d�e�e�e�f�l�G��H����V��L����u�d�d�d�f�l�F��I����V��_�D��e�d�e�y�]�}�W��H����W��_�E��e�d�d�d�f�l�G��I���F�^�E��e�e�e�e�g�m�G��H����W��^�W���u�u�w�e�g�m�G��I����V��_�D��d�d�e�d�u�}�W���[����V��^�E��e�e�e�e�f�l�F��I����FǻN��E��e�e�e�e�f�l�F��I����W��_�E��y�_�u�u�g�m�G��I����W��_�D��d�d�d�e�g�m�[�ԜY���V��^�E��e�e�d�e�f�l�F��H����V�d��U���e�e�e�e�g�l�F��I����W��_�D��d�w�u�u�w��G��I����W��_�D��e�d�d�d�f�m�F���Y���D��^�E��e�d�e�d�g�l�G��H����V��L����u�e�e�e�g�m�F��I����W��_�D��e�e�d�y�]�}�W��I����V��^�D��d�d�d�d�f�l�G��H���F�^�E��e�e�e�e�f�l�G��H����W��^�W���u�u�w�e�g�m�G��I����V��^�D��d�d�e�e�u�}�W���[����V��^�E��d�d�d�e�f�l�F��I����FǻN��E��e�e�e�d�g�m�F��H����W��_�E��y�_�u�u�g�m�G��I����V��_�E��d�d�d�e�g�l�[�ԜY���V��^�E��d�e�d�e�f�l�F��H����V�d��U���e�e�e�e�f�m�G��I����W��_�D��d�w�u�u�w��G��I����V��_�D��e�d�d�d�f�m�F���Y���D��^�E��e�e�d�d�f�l�G��H����V��L����u�e�e�e�g�m�G��H����W��_�D��e�e�e�y�]�}�W��I����V��_�D��d�e�d�d�f�l�G��H���F�^�E��e�d�d�e�g�m�F��H����W��^�W���u�u�w�e�g�m�G��H����W��^�D��d�d�e�d�u�}�W���[����V��_�D��d�e�d�e�f�l�F��I����FǻN��E��e�e�e�e�f�m�G��H����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�e�f�l�[�ԜY���V��^�D��d�e�e�e�f�l�F��H����W�d��U���e�e�e�e�f�m�F��H����W��_�D��d�w�u�u�w��G��I����V��^�D��d�d�d�d�f�m�F���Y���D��^�E��d�d�e�d�g�l�G��H����V��L����u�e�e�e�g�m�F��I����W��_�D��e�d�d�y�]�}�W��I����V��^�D��e�d�d�d�f�l�G��I���F�^�E��e�d�d�d�g�l�F��H����W��^�W���u�u�w�e�g�m�G��H����V��_�D��d�d�d�e�u�}�W���[����V��_�D��e�d�d�e�f�l�F��H����FǻN��E��e�e�e�d�f�l�G��H����W��_�E��y�_�u�u�g�m�G��H����V��^�E��d�d�d�e�f�m�[�ԜY���V��^�E��d�e�e�e�g�l�F��H����W�d��U���e�e�e�e�g�m�F��H����W��_�D��e�w�u�u�w��G��I����V��^�E��e�d�d�d�f�l�F���Y���D��^�E��e�d�d�d�f�m�G��H����W��L����u�e�e�e�g�l�G��I����W��_�D��d�e�e�y�]�}�W��I����W��_�E��d�e�d�d�f�l�F��H���F�^�E��e�e�d�e�g�m�G��H����W��^�W���u�u�w�e�g�m�G��H����W��_�D��d�d�e�d�u�}�W���[����V��^�E��e�d�d�d�f�l�F��I����FǻN��E��e�e�d�e�g�m�F��H����W��_�D��y�_�u�u�g�m�G��H����V��_�D��d�d�d�d�f�m�[�ԜY���V��^�E��d�e�d�e�g�l�F��H����V�d��U���e�e�e�e�g�l�F��I����W��_�D��e�w�u�u�w��G��I����W��^�D��e�d�d�d�f�l�F���Y���D��^�E��e�d�e�e�g�m�G��H����W��L����u�e�e�e�g�l�G��I����V��_�D��d�d�e�y�]�}�W��I����W��_�D��d�e�d�d�f�l�F��I���F�^�E��e�e�d�e�f�l�F��H����W��_�W���u�u�w�e�g�m�G��H����W��^�E��e�e�e�e�u�}�W���[����V��^�D��d�e�d�d�g�m�G��I����FǻN��E��e�e�d�e�f�m�G��H����V��^�E��y�_�u�u�g�m�G��H����V��_�D��e�e�e�e�f�m�[�ԜY���V��^�E��e�e�d�d�g�m�G��I����W�d��U���e�e�e�e�g�l�F��I����V��^�E��d�w�u�u�w��G��I����W��^�E��e�e�e�e�g�l�G���Y���D��^�E��e�e�e�e�f�l�G��I����W��L����u�e�e�e�g�l�G��I����W��^�E��e�e�e�y�]�}�W��I����W��^�E��e�d�e�e�g�m�G��I���F�^�E��e�e�d�e�f�m�G��I����V��_�W���u�u�w�e�g�m�G��I����V��^�E��e�e�d�d�u�}�W���[����V��^�D��e�d�d�e�g�m�G��I����FǻN��E��e�e�d�e�f�l�G��I����V��^�E��y�_�u�u�g�m�G��H����V��^�D��e�e�e�d�g�m�[�ԜY���V��^�E��d�e�d�e�f�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��d�e�e�e�g�m�F���Y���D��^�E��d�d�e�d�f�m�F��I����W��L����u�e�e�e�g�m�F��H����W��^�E��d�e�d�y�]�}�W��I����V��^�D��e�e�e�e�g�m�F��I���F�^�E��e�d�d�d�g�m�G��I����V��_�W���u�u�w�e�g�m�G��H����W��_�E��e�e�d�e�u�}�W���[����V��_�D��d�d�e�d�g�m�G��H����FǻN��E��e�e�e�d�f�m�F��I����V��^�D��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�D��e�e�e�d�g�m�G��I����V�d��U���e�e�e�e�f�l�F��I����V��^�D��d�w�u�u�w��G��I����W��_�D��d�e�e�e�f�m�G���Y���D��^�E��e�e�d�e�g�l�F��I����V��L����u�e�e�e�g�m�G��H����W��^�E��e�d�e�y�]�}�W��I����V��_�D��d�d�e�e�g�m�G��H���F�^�E��e�d�e�d�g�l�F��I����V��^�W���u�u�w�e�g�m�G��H����W��_�E��e�d�d�e�u�}�W���[����V��^�D��e�e�e�d�g�m�G��H����FǻN��E��e�e�e�d�g�m�F��H����V��_�E��y�_�u�u�g�m�G��I����W��_�D��e�e�e�e�f�m�[�ԜY���V��^�E��e�d�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�D��e�w�u�u�w��G��I����W��^�D��d�e�e�e�f�l�F���Y���D��^�E��e�d�e�e�g�m�G��I����W��L����u�e�e�e�g�m�G��H����W��^�E��d�e�e�y�]�}�W��I����V��_�E��e�d�e�e�g�m�F��I���F�^�E��e�e�e�d�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�d�e�d�u�}�W���[����W��_�D��d�e�e�e�g�m�G��I����FǻN��D��d�d�d�d�g�l�G��I����V��_�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�d�g�l�[�ԜY���W��_�D��d�e�e�e�g�m�G��I����W�d��U���d�d�d�d�f�m�G��I����V��^�D��e�w�u�u�w��F��H����W��_�D��e�e�e�e�f�m�G���Y���D��_�D��e�e�d�e�f�m�F��I����V��L����u�d�d�d�f�l�G��I����W��^�E��d�d�e�y�]�}�W��H����W��^�E��e�e�e�e�g�m�F��I���F�_�D��d�e�d�d�f�m�F��I����V��_�W���u�u�w�d�f�l�F��H����V��^�E��e�d�e�e�u�}�W���[����W��^�E��e�d�e�d�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��I����V��_�D��y�_�u�u�f�l�F��H����V��_�E��e�e�e�d�f�m�[�ԜY���W��_�E��d�e�d�e�g�m�G��I����V�d��U���d�d�d�d�g�l�G��H����V��^�D��e�w�u�u�w��F��H����W��_�D��e�e�e�e�f�m�F���Y���D��_�D��e�d�d�d�g�l�F��I����V��L����u�d�d�d�f�l�G��I����V��^�E��d�e�d�y�]�}�W��H����V��_�D��e�e�e�e�g�m�F��I���F�_�D��d�d�d�e�g�l�F��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�d�e�e�u�}�W���[����W��_�D��d�d�e�e�g�m�G��I����FǻN��D��d�d�e�d�g�l�F��I����V��_�E��y�_�u�u�f�l�F��I����V��^�D��e�e�e�e�f�l�[�ԜY���W��_�D��e�d�e�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�D��e�w�u�u�w��F��H����V��_�D��d�e�e�e�f�l�G���Y���D��_�D��e�d�d�d�g�m�G��I����W��L����u�d�d�d�f�m�G��I����W��^�E��e�e�e�y�]�}�W��H����V��^�E��d�d�e�e�g�m�G��H���F�_�D��d�e�d�e�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�d�e�d�u�}�W���[����W��^�E��d�e�d�e�g�m�G��I����FǻN��D��d�d�e�d�f�m�G��H����V��_�D��y�_�u�u�f�l�F��I����V��_�D��e�e�e�e�g�l�[�ԜY���W��_�E��d�e�e�d�g�m�G��I����W�d��U���d�d�d�d�g�m�G��I����V��^�D��e�w�u�u�w��F��H����W��^�E��d�e�e�e�g�l�F���Y���D��_�D��e�d�e�e�f�l�F��I����W��L����u�d�d�d�f�m�G��I����V��^�E��d�e�d�y�]�}�W��H����V��^�E��d�d�e�e�g�m�F��I���F�_�D��d�e�e�d�f�m�F��I����V��^�W���u�u�w�d�f�l�F��I����W��^�E��e�e�e�d�u�}�W���[����W��^�D��e�e�e�d�g�m�G��I����FǻN��D��d�d�e�e�g�l�F��H����V��^�E��y�_�u�u�f�l�F��I����V��^�D��e�e�e�d�g�l�[�ԜY���W��_�E��e�d�d�d�g�m�G��I����W�d��U���d�d�d�d�g�m�G��H����V��^�E��e�w�u�u�w��F��H����V��^�D��d�e�e�e�g�l�F���Y���D��_�D��d�d�d�d�g�m�G��I����W��L����u�d�d�d�f�l�F��H����V��^�E��e�d�d�y�]�}�W��H����W��_�E��d�e�e�e�g�m�G��H���F�_�D��e�d�d�d�f�l�F��I����V��^�W���u�u�w�d�f�l�G��H����W��^�E��e�e�e�e�u�}�W���[����W��_�D��d�d�d�e�f�l�F��H����FǻN��D��d�d�d�d�f�l�G��I����W��_�D��y�_�u�u�f�l�F��H����W��^�E��d�d�d�d�g�l�[�ԜY���W��_�E��e�e�e�e�f�l�F��H����V�d��U���d�d�d�d�g�m�G��I����W��_�D��d�w�u�u�w��F��H����V��^�D��e�d�d�d�f�m�G���Y���D��_�D��e�e�e�e�f�l�G��H����V��L����u�d�d�d�f�m�G��H����V��_�D��d�e�e�y�]�}�W��H����V��_�E��d�d�d�d�f�l�G��I���F�_�D��d�e�e�e�f�l�G��H����W��^�W���u�u�w�d�f�l�F��I����W��^�D��d�d�d�e�u�}�W���[����W��^�E��e�d�d�e�f�l�F��I����FǻN��D��d�d�e�e�g�m�F��I����W��_�D��y�_�u�u�f�l�F��I����V��^�D��d�d�d�e�g�l�[�ԜY���W��_�E��d�e�d�d�g�l�F��H����V�d��U���d�d�d�d�g�m�G��I����W��_�E��d�w�u�u�w��F��H����V��_�D��d�d�d�d�g�l�G���Y���D��_�D��d�d�e�d�f�m�G��H����W��L����u�d�d�d�f�m�F��H����W��_�D��d�e�e�y�]�}�W��H����V��^�E��e�d�d�d�f�l�F��I���F�_�D��d�e�d�e�f�l�F��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��d�e�e�d�u�}�W���[����W��_�E��d�d�d�e�f�l�F��I����FǻN��D��d�d�e�e�f�l�F��H����W��^�D��y�_�u�u�f�l�F��I����W��^�D��d�d�d�e�f�m�[�ԜY���W��_�D��e�d�d�d�g�l�F��H����V�d��U���d�d�d�d�f�m�G��H����W��_�E��e�w�u�u�w��F��H����V��_�E��d�d�d�d�g�m�F���Y���D��_�D��d�d�d�e�g�m�G��H����V��L����u�d�d�d�f�m�F��H����V��_�D��e�e�e�y�]�}�W��H����V��_�E��e�d�d�d�f�l�G��H���F�_�D��d�e�e�d�g�l�G��H����V��_�W���u�u�w�d�f�l�F��I����V��_�D��d�d�d�e�u�}�W���[����W��^�E��d�d�e�d�f�l�F��H����FǻN��D��d�d�d�d�g�m�G��I����W��_�E��y�_�u�u�f�l�F��H����V��_�E��d�d�e�d�g�l�[�ԜY���W��_�E��e�e�d�e�f�l�F��I����V�d��U���d�d�d�d�g�l�G��I����W��_�D��d�w�u�u�w��F��H����V��^�D��e�d�d�d�f�m�G���Y���D��_�D��e�d�d�e�f�l�G��H����V��L����u�d�d�d�f�l�G��I����V��_�D��d�e�d�y�]�}�W��H����W��^�D��e�e�d�d�f�m�F��I���F�_�D��d�d�e�e�f�l�F��H����V��^�W���u�u�w�d�f�l�F��H����W��^�D��d�d�e�e�u�}�W���[����V��^�E��e�e�e�e�f�l�F��H����FǻN��E��e�e�e�e�f�l�G��H����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�e�e�f�l�[�ԜY���V��^�E��d�e�d�d�f�l�F��I����W�d��U���e�e�e�e�g�m�G��H����W��_�D��e�w�u�u�w��G��I����W��_�D��d�d�d�d�f�l�G���Y���D��^�E��d�d�d�d�g�m�G��H����W��L����u�e�e�e�g�m�G��I����W��_�D��e�e�d�y�]�}�W��I����V��^�D��d�e�d�d�f�m�G��H���F�^�E��e�d�d�d�g�l�F��H����V��^�W���u�u�w�e�g�m�G��I����V��^�D��d�d�d�d�u�}�W���[����V��_�E��d�e�d�e�f�l�F��H����FǻN��E��e�e�e�d�f�l�G��H����W��_�E��y�_�u�u�g�m�G��H����V��^�D��d�d�e�e�g�l�[�ԜY���V��^�E��e�d�e�d�f�l�F��I����W�d��U���e�e�e�e�g�l�F��I����W��_�D��e�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�G���Y���D��^�E��d�e�d�d�f�l�F��H����W��L����u�e�e�e�g�l�F��I����W��_�D��e�d�e�y�]�}�W��I����W��^�D��e�d�d�d�f�m�G��I���F�^�E��e�d�d�e�f�m�G��H����V��_�W���u�u�w�e�g�m�G��H����W��^�D��d�d�e�e�u�}�W���[����V��_�E��e�e�e�d�f�l�F��I����FǻN��E��e�e�d�d�f�l�G��I����W��_�E��y�_�u�u�g�m�G��H����V��^�E��d�d�e�d�f�m�[�ԜY���V��^�E��e�d�d�d�g�l�F��I����W�d��U���e�e�e�d�g�m�G��I����W��_�D��d�w�u�u�w��G��I����W��^�D��e�d�d�d�f�l�G���Y���D��^�E��e�d�e�d�f�l�F��H����W��L����u�e�e�e�g�m�F��I����W��_�D��d�e�d�y�]�}�W��I����V��_�E��e�e�d�d�f�m�F��H���F�^�E��d�e�d�d�g�m�G��H����V��_�W���u�u�w�e�g�m�F��H����V��^�D��d�e�e�e�u�}�W���[����V��_�E��d�e�e�d�f�l�F��I����FǻN��E��e�e�e�e�f�m�G��I����W��^�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�e�f�l�[�ԜY���V��^�D��e�d�e�d�f�l�F��H����W�d��U���e�e�e�d�f�m�G��H����W��_�E��d�w�u�u�w��G��I����V��^�E��e�d�d�d�g�l�F���Y���D��^�E��d�d�d�e�g�l�G��H����V��L����u�e�e�e�g�m�F��H����W��_�D��d�e�d�y�]�}�W��I����V��_�D��e�e�d�d�f�l�F��H���F�^�E��d�d�d�d�g�m�G��H����W��^�W���u�u�w�e�g�m�F��I����V��^�D��d�e�d�d�u�}�W���[����V��^�E��d�d�e�e�f�l�F��H����FǻN��E��e�e�d�e�f�l�F��I����W��_�E��y�_�u�u�g�m�G��H����W��_�E��d�d�d�e�g�l�[�ԜY���V��^�E��e�d�e�e�f�l�F��H����V�d��U���e�e�e�d�g�l�F��I����W��_�D��e�w�u�u�w��G��I����W��^�D��e�d�d�d�f�l�G���Y���D��^�E��e�d�e�e�g�m�G��H����V��L����u�e�e�e�g�l�G��H����W��_�D��d�e�d�y�]�}�W��I����W��_�D��e�e�d�d�f�l�F��I���F�^�E��d�e�d�d�g�l�G��H����W��^�W���u�u�w�e�g�m�F��H����V��^�D��d�d�d�e�u�}�W���[����V��^�D��e�d�e�d�g�m�G��I����FǻN��E��e�e�d�e�f�m�F��H����V��^�E��y�_�u�u�g�m�G��H����W��_�D��e�e�e�e�f�l�[�ԜY���V��^�E��e�e�e�d�f�m�G��I����V�d��U���e�e�e�d�g�l�G��I����V��^�E��e�w�u�u�w��G��I����W��^�D��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�f�l�F��I����V��L����u�e�e�e�g�l�G��I����V��^�E��d�e�e�y�]�}�W��I����W��_�E��e�e�e�e�g�m�F��H���F�^�E��d�e�e�e�g�m�F��I����V��_�W���u�u�w�e�g�m�F��I����W��_�E��e�d�e�d�u�}�W���[����V��^�E��e�d�e�d�g�m�G��I����FǻN��E��e�e�e�d�f�m�G��I����V��_�E��y�_�u�u�g�m�G��I����W��_�D��e�e�e�e�f�l�[�ԜY���V��^�D��e�e�d�d�f�m�G��I����V�d��U���e�e�e�d�f�m�G��I����V��^�D��d�w�u�u�w��G��I����V��_�D��d�e�e�e�f�m�F���Y���D��^�E��e�d�d�d�f�l�F��I����W��L����u�e�e�e�g�m�G��I����W��^�E��d�d�e�y�]�}�W��I����V��_�E��d�e�e�e�g�l�G��H���F�^�E��d�d�e�e�f�m�F��I����W��_�W���u�u�w�e�g�m�F��H����V��^�E��e�e�e�d�u�}�W���[����V��^�E��e�e�e�e�g�m�G��H����FǻN��E��e�e�e�d�g�l�F��H����V��^�D��y�_�u�u�g�m�G��I����V��^�E��e�e�d�d�g�l�[�ԜY���V��^�E��e�d�e�e�f�m�G��H����V�d��U���e�e�e�d�g�m�G��I����V��^�E��d�w�u�u�w��G��I����W��^�D��d�e�e�e�g�l�F���Y���D��^�E��d�e�e�e�g�l�F��I����W��L����u�e�e�e�g�l�F��I����V��^�E��d�d�d�y�]�}�W��I����W��_�D��e�d�e�e�g�l�G��I���F�^�E��e�d�e�d�g�m�F��I����W��_�W���u�u�w�e�g�m�G��H����V��_�E��e�d�e�d�u�}�W���[����V��^�E��e�d�e�e�g�m�G��H����FǻN��E��e�e�d�d�g�m�F��I����V��_�D��y�_�u�u�g�m�G��H����W��_�E��e�e�d�e�f�m�[�ԜY���V��^�E��e�d�e�e�f�m�G��H����W�d��U���e�e�e�e�f�l�G��I����V��^�D��d�w�u�u�w��G��I����V��^�E��d�e�e�e�f�m�G���Y���D��^�E��e�d�e�e�g�m�F��I����V��L����u�e�e�e�g�m�G��H����V��^�E��d�e�e�y�]�}�W��I����V��_�E��d�e�e�e�g�l�F��I���F�^�E��e�e�e�d�f�l�F��I����W��_�W���u�u�w�e�g�m�G��H����W��_�E��e�d�d�e�u�}�W���[����V��^�D��d�d�d�e�g�m�G��H����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�e�g�l�[�ԜY���W��_�D��d�d�e�e�g�m�G��I����V�d��U���d�d�d�d�f�m�F��H����V��^�E��d�w�u�u�w��F��H����W��^�E��d�e�e�d�g�m�G���Y���D��_�D��d�d�d�e�g�l�F��I����V��L����u�d�d�d�f�l�G��I����V��^�E��e�d�d�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��_�W���u�u�w�d�f�l�F��I����V��_�E��d�e�e�e�u�}�W���[����W��_�D��e�e�e�d�g�m�F��I����FǻN��D��d�d�e�e�f�l�G��H����V��^�D��y�_�u�u�f�l�F��I����V��^�E��e�e�e�e�f�l�[�ԜY���W��_�E��e�d�e�d�g�m�G��I����W�d��U���d�d�d�d�g�l�G��I����V��^�E��e�w�u�u�w��F��H����V��^�E��e�e�e�d�g�m�F���Y���D��_�D��d�d�e�e�g�m�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�d�y�]�}�W��H����W��^�D��d�e�e�e�g�m�G��I���F�_�D��e�d�e�d�f�l�F��I����W��_�W���u�u�w�d�f�l�G��H����W��_�E��e�d�d�e�u�}�W���[����W��^�D��d�e�e�d�g�m�G��H����FǻN��D��d�d�d�e�f�m�F��I����V��_�E��y�_�u�u�f�l�F��H����W��_�D��e�e�d�d�g�m�[�ԜY���W��_�D��e�d�e�e�f�m�G��H����V�d��U���d�d�d�e�f�m�F��I����V��^�D��e�w�u�u�w��F��H����W��^�E��e�e�e�e�f�m�F���Y���D��_�D��e�e�e�d�f�l�G��I����V��L����u�d�d�d�f�m�G��H����V��^�E��e�d�d�y�]�}�W��H����V��^�D��d�d�e�e�g�l�G��I���F�_�D��e�e�e�e�g�l�F��I����W��^�W���u�u�w�d�f�l�G��H����W��_�E��e�d�e�e�u�}�W���[����W��^�E��e�d�e�e�g�m�G��I����FǻN��D��d�d�e�e�g�m�G��H����V��^�D��y�_�u�u�f�l�F��H����V��_�D��e�e�d�d�g�l�[�ԜY���W��^�D��d�d�d�d�g�m�G��H����V�d��U���d�d�d�d�f�m�G��H����V��^�E��e�w�u�u�w��F��H����W��_�E��d�e�e�e�g�m�G���Y���D��_�E��e�d�d�d�f�l�F��I����W��L����u�d�d�d�g�l�G��H����W��^�E��e�e�d�y�]�}�W��H����W��_�D��d�e�e�e�g�l�G��H���F�_�D��d�e�d�d�f�l�F��I����W��^�W���u�u�w�d�f�l�F��I����W��^�E��e�d�d�e�u�}�W���[����W��^�E��e�d�e�d�g�m�G��H����FǻN��D��d�e�d�d�g�m�F��H����V��_�D��y�_�u�u�f�l�F��H����W��_�E��e�e�e�d�g�m�[�ԜY���W��^�E��d�d�d�d�f�m�G��I����W�d��U���d�d�d�d�g�l�G��I����V��^�D��d�w�u�u�w��F��H����V��^�E��e�e�e�e�f�m�F���Y���D��_�E��e�d�e�d�f�l�F��I����W��L����u�d�d�d�g�l�G��I����W��^�E��d�e�e�y�]�}�W��H����W��^�D��e�d�e�e�g�m�F��H���F�_�D��d�e�e�e�f�l�F��I����V��_�W���u�u�w�d�f�l�F��I����W��^�E��e�e�d�e�u�}�W���[����W��_�D��d�e�e�d�g�m�G��I����FǻN��D��d�e�e�d�f�l�F��H����W��_�D��y�_�u�u�f�l�F��H����V��^�E��d�d�d�d�g�m�[�ԜY���W��^�E��e�e�e�d�g�l�F��H����W�d��U���d�d�d�d�g�m�F��H����W��_�D��d�w�u�u�w��F��H����V��_�E��d�d�d�d�f�l�F���Y���D��_�E��e�d�d�e�f�m�G��H����V��L����u�d�d�d�g�l�G��H����W��_�D��d�d�d�y�]�}�W��H����W��^�D��e�e�d�d�f�l�F��I���F�_�D��d�e�d�e�g�m�F��H����W��_�W���u�u�w�d�f�l�F��H����W��^�D��d�e�d�d�u�}�W���[����W��^�E��d�e�d�e�f�l�F��H����FǻN��D��d�e�d�d�f�m�F��H����W��^�D��y�_�u�u�f�l�F��H����V��^�D��d�d�e�d�f�l�[�ԜY���W��^�E��d�d�d�e�f�l�F��I����V�d��U���d�d�d�d�f�m�F��I����W��_�D��e�w�u�u�w��F��H����W��_�E��e�d�d�d�f�m�G���Y���D��_�E��e�d�d�d�f�l�F��H����W��L����u�d�d�d�g�l�F��H����V��_�D��e�d�d�y�]�}�W��H����W��^�D��d�d�d�d�f�m�G��I���F�_�D��d�d�d�d�f�l�F��H����V��^�W���u�u�w�d�f�l�G��I����V��_�D��d�e�e�d�u�}�W���[����W��^�D��e�e�e�e�f�l�F��I����FǻN��D��d�d�e�d�f�m�F��H����W��^�D��y�_�u�u�f�l�F��I����V��_�E��d�d�e�e�f�l�[�ԜY���W��_�D��e�e�d�e�g�l�F��I����W�d��U���d�d�d�e�f�l�G��I����W��_�D��d�w�u�u�w��F��H����V��_�E��e�d�d�e�f�l�F���Y���D��_�D��d�d�d�d�f�m�G��H����V��L����u�d�d�d�f�l�G��I����V��_�D��d�e�d�y�]�}�W��H����W��_�D��e�e�d�d�f�l�G��H���F�_�D��e�e�d�e�f�l�F��H����W��^�W���u�u�w�d�f�l�G��I����W��^�D��e�d�e�e�u�}�W���[����W��_�D��e�e�d�d�f�l�G��I����FǻN��D��d�d�d�d�f�m�F��I����W��^�D��y�_�u�u�f�l�F��I����W��^�D��d�d�d�d�g�l�[�ԜY���W��_�E��d�d�d�e�g�l�F��H����V�d��U���d�d�d�d�g�m�F��H����W��_�E��d�w�u�u�w��F��H����V��_�E��d�d�d�e�g�l�F���Y���D��_�D��e�d�e�d�f�l�F��H����W��L����u�d�d�d�f�m�F��I����W��_�D��e�e�e�y�]�}�W��H����W��^�D��d�e�d�d�f�l�G��H���F�_�D��d�e�d�d�f�l�G��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��e�e�e�d�u�}�W���[����W��_�D��e�d�e�e�f�l�G��I����FǻN��D��d�d�d�d�g�l�G��H����W��_�D��y�_�u�u�g�m�G��I����V��^�E��d�d�e�d�f�m�[�ԜY���V��^�E��e�e�e�d�g�l�F��I����V�d��U���e�e�e�e�g�l�G��I����W��_�D��e�w�u�u�w��G��I����V��^�D��e�d�d�e�f�m�F���Y���D��^�E��d�e�d�d�f�m�G��H����V��L����u�e�e�e�g�m�F��I����V��_�D��d�d�e�y�]�}�W��I����W��^�E��d�e�d�d�f�m�F��H���F�^�E��e�e�d�e�g�m�G��H����V��_�W���u�u�w�e�g�m�G��I����V��_�D��e�d�e�e�u�}�W���[����V��_�E��e�e�e�e�f�l�G��I����FǻN��E��e�e�d�d�f�m�F��H����W��_�D��y�_�u�u�g�m�G��I����W��^�E��d�d�e�d�f�m�[�ԜY���V��^�E��d�d�d�e�f�l�F��I����W�d��U���e�e�e�d�f�m�G��I����W��_�D��d�w�u�u�w��G��I����V��_�E��e�d�d�e�f�m�F���Y���D��^�E��d�d�d�d�f�m�G��H����W��L����u�e�e�e�g�l�G��H����W��_�D��d�e�d�y�]�}�W��I����W��_�E��e�d�d�d�f�m�F��H���F�^�E��d�d�e�d�g�l�F��H����V��_�W���u�u�w�e�g�m�F��H����V��_�D��e�d�d�d�u�}�W���[����V��_�E��d�d�d�e�f�l�G��I����FǻN��E��e�d�e�e�f�m�F��I����W��^�E��y�_�u�u�g�m�G��I����W��^�E��d�d�d�e�f�m�[�ԜY���V��_�E��e�e�e�d�g�l�F��H����W�d��U���e�e�e�e�f�l�G��I����W��_�E��e�w�u�u�w��G��I����V��_�E��d�d�d�e�g�l�F���Y���D��^�D��d�d�e�e�g�m�G��H����V��L����u�e�e�e�f�l�G��H����W��_�D��d�d�e�y�]�}�W��I����W��^�E��d�e�d�d�f�l�F��I���F�^�E��e�e�d�e�f�m�F��H����W��_�W���u�u�w�e�g�m�G��I����W��^�D��e�d�e�d�u�}�W���[����V��_�E��e�e�e�d�f�l�G��I����FǻN��E��e�d�d�d�g�m�F��H����W��_�D��y�_�u�u�g�m�G��I����W��_�D��d�d�d�d�g�l�[�ԜY���V��_�E��d�d�d�e�f�l�F��H����V�d��U���e�e�e�d�g�m�G��H����W��_�D��d�w�u�u�w��G��I����W��^�D��e�d�d�d�g�m�G���Y���D��^�D��e�e�d�d�f�m�G��H����V��L����u�e�e�e�f�m�G��H����V��_�D��e�d�e�y�]�}�W��I����V��^�E��d�d�d�d�f�m�F��H���F�^�E��d�d�d�e�f�m�G��H����V��^�W���u�u�w�e�g�m�F��H����W��_�D��d�e�d�d�u�}�W���[����V��^�D��d�d�d�e�f�l�F��I����FǻN��E��e�d�d�e�g�l�F��I����W��_�E��y�_�u�u�g�m�G��H����V��_�E��d�d�e�d�g�l�[�ԜY���V��_�E��d�e�d�e�g�l�F��I����V�N��X��>�:�3��:�/�E�ԜY���9l�T�����u��"�&��8��������g��z����o�<�!�2�%�g�W���Y���X*��R������1�-�:��4�:������F�d��U���i�>�:�0�#�2��������A2��D#��4���k�u�u�n�w�>�����Ƨ�Z��D�����;�0��'�?�.�6�������Z��P��O���u�u�x�i��:��������]��q�������!�k�w�}�E��Y���Z�������:�3��1�/�2�#���4����GV�N��N���6�;�!�;�w���������r
��T��'���c�!�o�u�]�}�W������U+��X����_�u�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�f�l�F��H����V��^�D��e�d�d�e�f�m�[�ԜY���W��^�E��d�d�d�d�f�m�G��H����W�d��U���d�d�e�e�f�l�G��I����V��_�D��d�w�u�u�w��F��I����V��_�E��d�e�e�e�g�l�F���Y���D��_�E��d�d�e�d�g�l�F��I����V��L����u�d�d�d�g�m�G��I����V��^�E��e�e�e�y�]�}�W��H����W��^�E��e�d�e�e�g�l�F��I���F�_�D��d�d�d�d�g�m�G��I����V��^�W���u�u�w�d�f�l�F��I����V��_�E��d�d�e�e�u�}�W���[����W��^�D��e�e�e�d�g�m�F��H����FǻN��D��e�d�d�d�f�m�G��I����V��_�E��y�_�u�u�f�l�G��H����V��^�D��e�e�d�e�g�l�[�ԜY���W��_�E��e�d�e�e�f�m�G��H����W�d��U���d�d�d�d�g�m�G��H����V��^�D��d�w�u�u�w��F��H����V��^�D��d�e�e�e�f�m�F���Y���D��_�D��e�e�e�d�g�m�G��I����V��L����u�d�d�e�f�l�G��I����V��^�E��e�e�d�y�]�}�W��H����W��^�E��d�e�d�d�f�l�G��H���F�_�D��d�e�e�e�g�l�G��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�e�d�e�u�}�W���[����W��^�D��d�d�d�e�f�l�F��H����FǻN��D��e�d�d�d�g�m�F��H����W��_�D��y�_�u�u�f�l�G��H����V��^�D��d�d�e�d�f�m�[�ԜY���W��_�E��d�d�d�d�g�l�F��I����W�d��U���d�d�d�d�f�m�F��H����W��_�D��d�w�u�u�w��F��H����V��_�E��e�d�d�e�f�m�G���Y���D��_�D��d�e�e�d�g�m�G��H����V��L����u�d�d�d�g�m�G��I����W��_�D��d�d�d�y�]�}�W��H����V��^�E��e�d�d�d�f�l�G��H���F�_�D��e�e�d�e�g�m�F��H����W��^�W���u�u�w�d�f�m�G��H����W��_�D��e�d�e�e�u�}�W���[����V��_�D��d�d�d�e�f�l�G��H����FǻN��D��d�e�d�e�f�m�F��H����W��_�E��y�_�u�u�f�l�F��H����V��_�E��d�d�e�d�f�l�[�ԜY���W��^�D��d�e�e�e�g�l�F��I����V�d��U���d�d�e�e�f�m�G��H����W��_�E��e�w�u�u�w��F��I����V��_�E��e�d�d�d�f�l�F���Y���D��_�E��d�e�e�e�g�m�F��H����V��L����u�d�d�d�g�m�G��H����W��_�E��e�d�d�y�]�}�W��H����V��_�D��d�e�d�d�g�l�G��H���F�_�D��d�e�e�d�f�m�F��H����W��^�W���u�u�w�d�f�m�F��H����W��_�D��d�e�d�d�u�}�W���[����V��_�E��d�e�e�e�f�l�F��H����FǻN��D��d�e�d�d�f�m�G��I����W��^�D��y�_�u�u�f�l�F��I����W��_�E��d�e�d�d�g�l�[�ԜY���W��_�D��e�e�e�e�g�l�F��H����W�d��U���d�d�e�e�f�m�F��H����W��^�E��d�w�u�u�w��F��I����W��^�E��d�d�d�d�g�m�F���Y���D��_�D��d�d�e�d�f�m�G��H����V��L����u�d�d�d�f�l�F��I����V��_�E��e�e�d�y�]�}�W��H����V��_�D��e�e�d�d�g�l�G��I���F�_�D��d�e�d�d�g�l�G��H����W��^�W���u�u�w�d�f�m�F��H����W��^�D��d�e�e�e�u�}�W���[����V��^�E��d�e�d�e�f�l�F��I����FǻN��D��d�d�d�d�f�m�F��H����W��^�E��y�_�u�u�f�l�F��H����V��^�E��d�e�d�e�g�l�[�ԜY���W��_�D��d�e�d�d�f�l�F��H����V�d��U���d�d�d�e�g�m�G��H����W��^�E��d�w�u�u�w��F��H����V��_�D��d�d�d�d�g�m�G���Y���D��_�E��d�e�d�d�g�m�F��H����V��L����u�d�d�d�g�l�G��I����V��_�E��e�e�d�y�]�}�W��H����W��^�E��e�e�d�d�g�l�G��H���F�_�D��e�d�e�d�g�l�G��H����W��_�W���u�u�w�d�f�l�F��I����W��_�D��d�e�e�e�u�}�W���[����W��^�E��d�e�d�e�f�l�F��I����FǻN��D��d�e�e�e�g�l�F��H����W��^�E��y�_�u�u�f�l�F��I����W��_�E��d�e�d�d�g�l�[�ԜY���W��^�E��d�d�e�e�g�l�F��H����W�d��U���d�d�d�d�f�m�G��I����W��^�D��d�w�u�u�w��F��H����V��^�D��e�d�d�d�f�l�G���Y���D��_�D��e�d�e�d�g�l�F��H����W��L����u�d�d�d�f�m�F��H����W��_�E��d�e�d�y�]�}�W��H����V��_�D��d�e�d�d�g�l�F��I���F�_�D��e�d�e�d�g�l�F��H����W��^�W���u�u�w�d�f�l�G��I����W��_�D��e�e�e�e�u�}�W���[����W��^�D��d�e�d�e�f�l�G��I����FǻN��D��d�d�d�e�f�l�G��I����W��^�E��y�_�u�u�f�l�F��H����V��^�D��d�d�e�d�g�l�[�ԜY���W��_�E��d�d�d�d�g�l�F��I����V�d��U���d�d�d�d�g�m�G��H����W��_�E��e�w�u�u�w��F��H����W��_�E��d�d�d�e�f�m�F���Y���D��_�D��e�d�e�d�g�l�G��H����W��L����u�d�d�d�f�m�F��H����V��_�D��e�d�e�y�]�}�W��H����W��_�E��e�e�d�d�f�m�F��I���F�_�D��d�e�e�d�g�l�F��H����V��^�W���u�u�w�d�f�l�F��H����W��_�D��e�e�e�e�u�}�W���[����W��_�E��e�e�d�d�f�l�G��I����FǻN��D��d�d�d�d�f�l�F��I����W��^�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�g�l�[�ԜY���V��^�E��d�e�d�d�f�l�F��H����W�d��U���e�e�e�e�g�m�G��I����W��_�D��e�w�u�u�w��G��I����W��^�E��d�d�d�e�f�m�F���Y���D��^�E��e�d�d�d�g�m�F��H����W��L����u�e�e�e�g�m�F��I����W��_�D��d�e�e�y�]�}�W��I����V��^�D��e�e�d�d�f�l�F��I���F�^�E��e�e�e�e�f�m�F��H����W��_�W���u�u�w�e�g�m�G��H����V��^�D��d�e�e�e�u�}�W���[����V��^�D��d�d�e�d�f�l�F��H����FǻN��E��e�e�d�d�f�m�F��H����W��^�E��y�_�u�u�g�m�G��H����W��^�D��d�d�e�d�f�m�[�ԜY���V��^�D��d�d�e�d�g�l�F��I����V�d��U���e�e�e�e�f�l�G��H����W��_�D��d�w�u�u�w��G��I����W��^�D��d�d�d�d�f�m�F���Y���D��^�E��d�d�e�d�g�l�G��H����W��L����u�e�e�e�g�l�F��H����W��_�D��d�e�e�y�]�}�W��I����W��_�D��d�e�d�d�f�m�F��I���F�^�E��d�e�e�e�f�l�F��H����V��_�W���u�u�w�e�g�m�F��I����V��^�D��d�e�e�d�u�}�W���[����V��^�E��d�d�d�d�f�l�F��I����FǻN��E��e�e�e�e�f�m�G��I����W��^�D��y�_�u�u�g�m�G��I����W��^�E��d�d�d�d�g�l�[�ԜY���V��^�E��d�e�d�d�f�l�F��H����V�d��U���e�e�e�d�g�m�G��I����W��_�E��d�w�u�u�w��G��I����V��_�D��d�d�d�d�g�l�F���Y���D��^�E��d�e�e�d�f�m�F��H����V��L����u�e�e�e�g�m�F��H����V��_�D��e�e�e�y�]�}�W��I����V��^�E��e�d�d�d�f�l�G��I���F�^�E��d�e�d�e�g�l�G��H����W��^�W���u�u�w�e�g�m�F��H����W��_�D��d�d�e�e�u�}�W���[����V��^�D��d�d�e�d�f�l�F��I����FǻN��E��e�e�e�d�f�l�F��I����W��_�E��y�_�u�u�g�m�G��I����W��_�D��d�d�d�d�f�l�[�ԜY���V��^�E��e�d�d�e�f�m�G��I����V�d��U���e�e�e�d�g�l�G��H����V��^�E��e�w�u�u�w��G��I����W��_�D��e�e�e�e�g�l�G���Y���D��^�E��d�d�e�e�g�m�F��I����W��L����u�e�e�e�g�m�F��H����W��^�E��e�d�e�y�]�}�W��I����V��^�E��d�e�e�e�g�m�F��H���F�^�E��d�e�d�e�g�m�G��I����V��^�W���u�u�w�e�g�m�F��I����W��^�E��e�e�e�d�u�}�W���[����V��^�D��e�d�e�d�g�m�G��H����FǻN��E��e�e�e�d�f�m�F��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�d�f�l�[�ԜY���V��^�E��e�d�d�d�f�m�G��I����W�d��U���e�e�e�d�g�l�F��H����V��^�D��e�w�u�u�w��G��I����W��_�D��d�e�e�e�f�m�F���Y���D��^�E��e�e�e�d�f�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�d�d�y�]�}�W��I����V��_�D��e�d�e�e�g�m�G��H���F�^�E��d�e�e�d�g�m�F��I����V��^�W���u�u�w�e�g�m�F��I����V��^�E��e�d�d�e�u�}�W���[����V��_�D��d�e�e�e�g�m�G��H����FǻN��E��e�e�d�d�g�l�G��H����V��_�E��y�_�u�u�g�m�G��H����V��^�D��e�e�e�e�f�m�[�ԜY���V��^�D��e�d�d�e�f�m�G��I����W�d��U���e�e�e�e�f�m�F��I����V��^�D��e�w�u�u�w��G��I����W��_�E��d�e�e�e�f�l�F���Y���D��^�E��e�d�d�e�g�m�F��I����W��L����u�e�e�e�g�l�G��I����W��^�E��e�d�d�y�]�}�W��I����W��_�E��e�d�e�e�g�m�G��H���F�^�E��e�d�e�e�g�l�F��I����V��_�W���u�u�w�e�g�m�G��I����W��_�E��e�d�e�e�u�}�W���[����V��^�D��e�d�e�d�g�m�G��I����FǻN��E��e�e�d�d�g�l�G��H����V��_�E��y�_�u�u�g�m�G��H����V��^�D��e�e�e�d�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�F��I����V��^�D��d�w�u�u�w��G��I����W��^�D��d�e�e�e�f�l�F���Y���D��^�E��e�d�e�e�g�m�F��I����W��L����u�e�e�e�g�l�G��H����W��^�E��e�d�e�y�]�}�W��I����W��_�D��d�e�e�e�g�m�G��I���F�^�E��e�e�e�d�f�l�F��I����V��_�W���u�u�w�e�g�m�G��I����W��_�E��e�d�d�e�u�}�W���[����V��_�D��d�e�d�e�g�m�G��H����FǻN��E��e�e�e�d�g�l�G��I����V��_�E��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�g�l�[�ԜY���V��^�D��d�e�d�d�g�m�G��I����V�d��U���e�e�e�e�f�m�F��I����V��^�D��e�w�u�u�w��G��I����V��^�D��e�e�e�e�f�l�G���Y���D��^�E��e�d�e�d�f�l�F��I����W��L����u�e�e�e�g�m�G��I����V��^�E��e�d�d�y�]�}�W��I����V��^�E��d�d�e�e�g�m�G��I���F�^�E��e�d�e�d�f�l�F��I����V��_�W���u�u�w�e�g�m�G��I����W��^�E��e�d�e�e�u�}�W���[����V��_�E��d�e�d�e�g�m�G��I����FǻN��E��e�e�e�e�g�l�G��H����V��_�E��y�_�u�u�g�m�G��I����W��^�D��e�e�e�e�g�l�[�ԜY���V��^�E��e�e�e�e�f�m�G��I����V�d��U���e�e�e�e�g�l�F��I����V��^�E��d�w�u�u�w��G��I����W��^�E��e�e�e�e�g�l�F���Y���D��^�E��d�d�d�d�g�l�G��I����W��L����u�e�e�e�g�m�F��H����W��^�E��d�d�e�y�]�}�W��I����V��^�D��d�d�e�e�g�m�F��H���F�^�E��e�e�e�d�g�l�G��I����V��^�W���u�u�w�e�g�m�G��I����V��_�E��e�e�d�d�u�}�W���[����V��^�D��e�e�d�e�g�m�G��H����FǻN��E��e�e�e�e�f�l�G��H����V��^�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�d�f�l�[�ԜY���V��^�E��d�d�e�d�g�m�G��I����V�d��U���e�e�e�e�g�l�G��H����V��^�E��e�w�u�u�w��G��I����W��^�E��d�e�e�e�g�m�G���Y���D��^�E��e�d�d�e�f�l�G��I����V��L����u�e�e�e�g�m�G��H����W��^�E��d�e�e�y�]�}�W��I����V��_�D��e�e�e�e�g�m�F��H���F�^�E��e�e�e�d�f�l�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�d�u�}�W���[����V��^�E��e�e�d�e�g�m�G��H����FǻN��E��e�e�e�e�g�l�G��H����V��^�D��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�f�l�[�ԜY���W��_�D��d�d�d�e�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��d�w�u�u�w��F��H����W��^�E��d�e�e�e�g�l�F���Y���D��_�D��d�d�d�e�g�m�F��I����W��L����u�d�d�d�f�l�F��H����V��^�E��e�e�d�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�d�d�e�g�m�F��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�d�u�}�W���[����W��_�E��d�e�e�e�g�m�G��I����FǻN��D��d�d�d�d�g�m�F��H����V��^�D��y�_�u�u�f�l�F��H����V��_�D��e�e�e�e�f�l�[�ԜY���W��_�D��d�e�e�d�g�m�G��I����W�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�G���Y���D��_�D��d�e�d�e�f�m�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��e�e�d�y�]�}�W��H����W��^�E��d�e�e�e�g�m�G��I���F�_�D��d�d�d�e�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����V��_�E��e�e�e�e�u�}�W���[����W��_�E��e�e�e�d�g�m�G��I����FǻN��D��d�d�d�d�g�l�G��I����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��e�d�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�G��I����V��^�E��e�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�F���Y���D��_�D��d�e�d�e�f�m�G��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�d�y�]�}�W��H����W��^�E��e�e�d�d�f�l�F��H���F�_�D��d�d�d�e�g�m�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�E��e�d�d�e�f�l�F��H����FǻN��D��d�d�d�d�g�l�G��H����W��_�D��y�_�u�u�f�l�F��H����W��_�E��d�d�d�d�f�m�[�ԜY���W��_�D��e�d�d�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��H����W��_�D��d�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�G���Y���D��_�D��d�e�e�d�f�m�F��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�d�y�]�}�W��H����W��^�D��e�e�d�d�f�l�F��H���F�_�D��d�d�d�d�f�l�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�e�u�}�W���[����W��_�E��d�d�e�d�f�l�F��H����FǻN��D��d�d�d�d�g�l�G��H����W��_�D��y�_�u�u�f�l�F��H����W��_�E��d�d�d�d�f�l�[�ԜY���W��_�D��d�d�d�e�g�l�F��H����W�d��U���d�d�d�d�f�l�G��I����W��_�D��e�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�G���Y���D��_�D��d�d�e�d�g�l�F��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�d�d�y�]�}�W��H����W��_�D��e�d�d�d�f�l�F��H���F�_�D��d�d�d�e�f�l�G��H����W��_�W���u�u�w�d�f�l�F��H����V��^�D��d�d�d�e�u�}�W���[����W��_�D��d�e�d�e�f�l�F��H����FǻN��D��d�d�d�d�f�l�F��H����W��_�D��y�_�u�u�f�l�F��H����W��_�D��d�d�d�d�f�m�[�ԜY���W��_�D��e�d�d�d�g�l�F��H����V�d��U���d�d�d�d�f�l�G��H����W��_�D��d�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�e�e�g�m�F��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�e�y�]�}�W��H����W��_�E��d�e�d�d�f�l�F��I���F�_�D��d�d�d�d�f�m�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�D��d�e�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�F��I����W��_�D��y�_�u�u�f�l�F��H����V��_�E��d�d�d�d�f�m�[�ԜY���W��_�D��d�e�e�e�f�l�F��H����V�d��U���d�d�d�d�f�l�F��H����W��_�D��d�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�F���Y���Z��t�����:�,�9�e�]�}�W��Y���F��Y������"�&��2�;����?����Z��T/��D��<�!�2�'�m�}�W���T�ڧ�\��C-�����1�-�:��>�����H���F��d��U���i�>�:�0�#�2��������A2��D#��4���k�u�u�n�w�>�����Ƨ�Z��D�����;�0��'�?�.�6�������Z��P��O���u�u�x�i��:��������]��q�������!�k�w�}�B��Y���Z�������:�3��1�/�2�#���4����GW�N��N���u�6�;�!�9�}�4�������A��C_��U����c�!�o�w�W�W���Tύ��V ��R�����d�_�u�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���V��^�E��e�e�e�e�g�m�G��I����V��B��U���w�e�e�e�g�m�G��I����V��^�E��e�e�w�u�w�}�U��I����V��^�E��e�e�e�e�g�m�G��[��ƹF�^�E��e�e�e�e�g�m�G��I����V��^�Y�ߊu�u�e�e�g�m�G��I����V��^�E��e�e�e�e�{�W�W���I����V��^�E��e�e�e�e�g�m�G��I���l�N��E��e�e�e�e�g�m�G��I����V��^�E���u�u�u�w�g�m�G��I����V��^�E��e�e�e�e�g��W���Y����V��^�E��e�e�e�e�g�m�G��I����D�=N��U��e�e�e�e�g�m�G��I����V��^�E��e�y�_�u�w�m�G��I����V��^�E��e�e�e�e�g�m�G��s���W��_�E��d�d�d�d�f�l�F��I����W��B��U���w�d�d�e�g�l�G��H����W��_�D��e�d�w�u�w�}�U��H����W��_�D��e�d�d�d�f�m�F��[��ƹF�_�D��e�e�d�e�f�l�G��H����V��^�Y�ߊu�u�d�d�f�m�G��I����W��^�D��d�e�d�d�{�W�W���H����V��^�D��d�e�d�d�f�m�F��I���l�N��D��e�d�d�e�g�m�G��I����V��^�D���u�u�u�w�f�l�G��H����W��^�E��d�e�e�e�g��W���Y����W��^�E��e�d�e�e�f�l�G��H����D�=N��U��d�d�d�d�g�m�G��I����W��_�D��e�y�_�u�w�l�F��H����W��^�E��d�d�d�d�g�m�G��s���W��_�D��d�e�e�e�g�m�F��H����V��B��U���w�d�d�e�f�l�G��H����W��_�D��e�d�w�u�w�}�U��H����V��^�D��e�e�d�e�g�l�F��[��ƹF�_�D��e�e�e�e�g�l�F��H����V��^�Y�ߊu�u�d�d�f�m�G��H����V��_�D��e�e�d�d�{�W�W���H����V��^�E��e�e�d�d�f�l�G��I���l�N��D��d�d�e�e�g�m�G��H����V��_�E���u�u�u�w�f�l�F��I����W��_�E��e�d�e�e�f��W���Y����W��_�D��e�d�d�d�f�l�G��H����D�=N��U��d�d�d�e�f�m�G��H����W��_�D��e�y�_�u�w�l�F��H����V��^�D��d�d�e�d�f�l�G��s���W��_�D��e�e�e�d�f�l�F��I����W��B��U���w�d�d�d�f�l�G��I����V��_�E��e�e�w�u�w�}�U��I����V��_�D��d�e�d�e�g�l�G��[��ƹF�^�E��d�d�d�e�g�l�G��H����V��^�Y�ߊu�u�e�e�g�m�G��I����V��_�E��d�e�d�d�{�W�W���I����V��^�D��d�e�d�d�g�l�F��I���l�N��E��e�e�d�d�g�l�F��I����W��^�E���u�u�u�w�g�m�G��H����V��^�D��d�d�e�d�f��W���Y����V��_�D��d�e�e�d�f�l�F��H����D�=N��U��e�e�e�e�g�m�F��I����W��^�D��e�y�_�u�w�m�G��I����V��_�E��d�e�d�e�f�l�F��s���V��^�D��d�d�d�d�g�l�F��H����V��B��U���w�e�e�d�f�l�F��H����W��^�D��d�d�w�u�w�}�U��I����V��^�E��d�d�d�d�f�l�G��[��ƹF�^�E��e�d�d�e�g�m�G��H����V��_�Y�ߊu�u�e�e�g�l�F��I����V��_�E��e�e�d�e�{�W�W���I����V��^�E��d�e�e�d�g�m�G��I���l�N��E��e�d�e�d�g�l�F��H����V��_�D���u�u�u�w�g�m�G��H����V��^�D��d�e�e�d�g��W���Y����V��^�E��d�e�e�e�f�l�F��I����D�=N��U��e�d�d�e�g�l�G��I����W��^�E��e�y�_�u�w�m�G��I����V��_�D��d�e�e�e�f�m�F��s���V��_�E��d�d�d�e�f�m�F��H����V��B��U���w�e�e�d�f�m�F��H����W��^�D��e�d�w�u�w�}�U��I����W��^�E��e�d�d�e�f�m�F��[��ƹF�^�D��e�d�d�d�g�l�G��H����W��^�Y�ߊu�u�e�e�f�l�F��I����V��_�E��e�d�d�d�{�W�W���I����V��^�D��d�d�d�d�g�l�G��I���l�N��E��e�d�e�d�f�l�G��H����W��_�D���u�u�u�w�g�l�G��H����W��_�D��e�e�d�e�f��W���Y����W��_�E��e�e�d�e�f�l�G��I����D�=N��U��e�e�e�e�g�l�G��I����W��^�D��d�y�_�u�w�m�G��I����V��^�D��d�e�d�e�g�l�G��s���V��^�D��d�e�e�d�g�m�F��H����V��B��U���w�e�d�d�g�m�G��H����W��^�E��d�e�w�u�w�}�U��H����V��_�D��e�e�d�e�f�l�F��[��ƹF�^�D��e�d�e�d�g�m�F��H����W��_�Y�ߊu�u�e�e�f�m�G��I����V��_�E��d�e�e�e�{�W�W���I����W��_�E��e�d�e�d�g�m�F��H���l�N��E��e�d�e�e�g�l�F��I����V��^�D���u�u�u�w�g�l�F��I����V��^�D��e�d�e�e�g��W���Y����W��^�D��d�e�e�e�g�l�G��H����D�=N��U��e�d�e�d�g�l�G��I����W��_�E��e�y�_�u�w�m�G��H����W��_�E��d�e�e�e�g�l�G��s���V��_�D��d�d�e�d�f�l�F��I����W��B��U���w�e�e�e�g�m�G��H����W��^�D��d�d�w�u�w�}�U��I����V��_�D��d�d�d�e�f�m�G��[��ƹF�^�E��e�d�d�e�f�l�F��H����V��_�Y�ߊu�u�e�d�g�l�G��H����W��^�E��e�d�e�e�{�W�W���I����V��^�E��d�d�d�d�g�m�G��H���l�N��E��d�d�d�e�f�l�G��I����V��^�D���u�u�u�w�g�m�F��I����W��^�D��e�d�e�d�f��W���Y����V��_�D��d�e�e�e�g�l�G��I����D�=N��U��d�d�e�e�g�m�G��H����W��_�D��e�y�_�u�w�m�F��I����W��_�E��d�e�e�e�f�m�G��s���V��_�D��e�e�e�d�f�m�F��I����W��B��U���w�e�e�e�g�l�F��H����V��^�D��e�d�w�u�w�}�U��I����W��^�D��d�d�d�e�f�l�F��[��ƹF�^�D��d�d�d�d�g�m�G��H����W��_�Y�ߊu�u�e�d�f�m�F��I����V��^�E��e�d�d�e�{�W�W���I����W��_�E��d�d�d�d�g�m�F��H���l�N��E��d�d�d�d�f�l�F��H����V��_�D���u�u�u�w�g�l�G��H����W��_�E��e�d�d�e�g��W���Y����W��_�D��e�d�d�d�g�l�G��H����D�=N��U��d�e�d�e�g�m�F��I����W��_�D��d�y�_�u�w�m�F��H����V��^�D��d�e�d�e�g�l�G��s���V��^�D��e�e�e�d�f�l�F��H����W��B��U���w�e�d�d�g�m�F��I����V��^�E��e�d�w�u�w�}�U��H����W��^�D��e�d�d�e�g�m�G��[��ƹF�^�E��e�e�e�d�g�m�G��H����V��_�Y�ߊu�u�e�d�g�l�G��H����V��_�E��d�d�e�e�{�W�W���I����W��_�D��e�e�e�d�g�l�G��H���l�N��E��e�e�e�d�g�l�G��H����W��_�D���u�u�u�w�g�l�G��H����V��^�E��e�d�d�d�g��W���Y����W��^�E��d�d�e�d�g�l�G��I����D�=N��U��d�d�d�e�g�m�G��H����W��_�E��d�y�_�u�w�m�F��H����V��_�D��d�e�e�e�g�m�F��s���V��_�E��d�d�d�e�g�m�F��I����W��B��U���w�e�d�d�f�m�F��I����W��^�E��e�e�w�u�w�}�U��H����W��^�E��d�d�d�d�g�l�G��[��ƹF�^�D��d�e�d�e�f�l�F��H����V��_�Y�ߊu�u�e�d�f�l�G��I����W��_�E��e�e�d�e�{�W�W���I����W��_�D��d�e�d�d�g�m�F��H���l�N��D��e�e�e�e�f�l�G��H����V��^�E���u�u�u�w�f�m�G��I����V��^�D��d�e�e�d�g��W���Y����V��_�E��e�e�d�d�f�l�F��H����D�=N��U��e�e�d�e�g�l�G��I����W��^�D��d�y�_�u�w�m�G��H����W��^�D��d�e�d�d�f�l�G��s���V��^�D��d�e�d�d�f�m�F��H����V��B��U���w�d�e�d�g�m�G��I����V��^�D��d�d�w�u�w�}�U��I����V��^�E��d�d�d�d�f�l�G��[��ƹF�_�E��d�d�d�d�f�l�G��H����V��_�Y�ߊu�u�e�e�g�m�G��I����V��^�D��d�e�d�d�{�W�W���I����V��_�E��d�d�d�d�f�m�F��H���l�N��D��d�e�d�d�f�l�G��H����V��_�D���u�u�u�w�f�m�F��I����V��_�D��e�d�e�e�f��W���Y����V��_�E��d�e�e�d�g�l�G��H����D�=N��U��e�e�d�e�f�l�F��I����W��^�D��d�y�_�u�w�m�G��H����V��_�D��d�d�d�d�g�l�G��s���V��_�E��e�e�d�e�g�l�F��H����V��B��U���w�d�e�e�g�l�G��I����W��_�D��e�d�w�u�w�}�U��I����V��^�D��e�e�d�e�f�m�G��[��ƹF�_�D��d�d�e�e�g�m�F��H����V��^�Y�ߊu�u�e�e�f�m�G��H����V��^�D��e�d�d�e�{�W�W���I����V��^�D��d�e�e�d�f�m�F��H���l�N��D��e�d�e�e�g�l�F��I����V��_�D���u�u�u�w�f�m�G��I����W��_�D��d�d�e�e�g��W���Y����V��_�E��e�e�e�e�g�l�F��H����D�=N��U��e�d�e�d�f�m�G��H����W��^�E��e�y�_�u�w�m�G��H����V��_�D��d�d�d�d�f�l�F��s���V��_�E��d�d�d�e�f�m�F��H����W��B��U���w�d�e�e�g�m�F��I����W��_�D��e�d�w�u�w�}�U��I����V��^�E��e�e�d�d�f�l�F��[��ƹF�_�D��e�e�d�d�g�m�G��I����V��^�Y�ߊu�u�e�e�f�l�G��I����V��_�E��d�e�e�d�{�W�W���I����W��^�D��d�d�d�e�g�m�F��I���l�N��D��e�d�d�d�g�m�F��H����V��^�D���u�u�u�w�f�m�G��H����W��^�E��e�d�e�d�g��W���Y����V��_�D��d�e�d�d�f�m�G��I����D�=N��U��e�d�e�d�g�l�F��H����V��^�D��e�y�_�u�w�m�G��I����W��^�E��e�e�d�d�g�l�F��s���V��_�D��e�e�e�d�f�l�G��H����W��B��U���w�d�e�e�g�l�F��H����V��^�D��d�e�w�u�w�}�U��I����V��^�D��e�e�e�e�f�l�F��[��ƹF�_�D��e�d�d�e�f�l�G��I����W��_�Y�ߊu�u�e�e�f�m�G��I����W��^�E��d�d�e�d�{�W�W���I����W��^�E��d�d�e�e�g�m�G��H���l�N��D��d�d�d�d�g�m�F��I����V��_�E���u�u�u�w�f�m�F��I����V��_�E��d�d�d�e�g��W���Y����V��^�D��e�e�e�d�f�m�F��I����D�=N��U��e�e�d�e�g�m�G��I����V��^�D��e�y�_�u�w�m�G��I����W��^�D��e�e�d�d�g�l�G��s���V��^�D��d�d�e�d�g�l�G��H����V��B��U���w�d�e�d�g�l�F��I����V��^�D��d�d�w�u�w�}�U��I����V��^�E��d�d�e�d�f�l�G��[��ƹF�_�E��e�e�e�e�f�m�G��I����V��_�Y�ߊu�u�e�e�g�l�G��H����V��^�D��e�d�d�e�{�W�W���I����W��_�D��e�d�d�e�f�m�F��H���l�N��D��e�e�d�d�f�l�G��H����V��^�E���u�u�u�w�f�m�G��H����V��_�D��e�d�d�d�f��W���Y����V��_�D��d�e�e�e�f�m�G��I����D�=N��U��e�e�e�d�g�l�F��H����V��_�D��e�y�_�u�w�m�F��H����W��_�E��e�d�d�e�f�m�G��s���V��_�D��e�d�d�d�f�l�G��H����V��B��U���w�e�d�d�g�m�F��H����W��_�E��d�e�w�u�w�}�U��H����W��^�E��d�d�e�e�g�l�F��[��ƹF�^�D��e�d�e�d�f�l�G��I����V��^�Y�ߊu�u�e�d�f�m�G��H����W��_�D��e�d�d�e�{�W�W���I����W��^�E��d�d�d�e�f�l�F��I���l�N��E��e�d�e�e�f�m�F��H����W��_�D���u�u�u�w�g�l�G��H����V��^�E��d�e�e�e�f��W���Y����W��_�D��e�d�e�e�g�m�F��H����D�=N��U��d�d�e�d�f�m�F��H����V��^�E��e�y�_�u�w�m�F��H����V��_�E��e�d�e�d�g�m�F��s���V��^�D��d�e�e�d�f�l�G��I����V��B��U���w�e�d�d�g�l�G��I����W��_�D��e�e�w�u�w�}�U��H����W��^�D��e�d�e�d�f�l�G��[��ƹF�^�E��d�e�d�d�g�m�G��I����W��_�Y�ߊu�u�e�d�g�l�F��I����W��^�D��d�e�d�e�{�W�W���I����W��_�D��d�d�d�e�f�m�F��I���l�N��E��e�e�e�e�f�m�G��H����V��_�D���u�u�u�w�g�l�G��I����W��_�E��d�e�e�e�f��W���Y����W��^�E��d�e�d�d�g�m�F��I����D�=N��U��d�d�d�e�g�l�F��H����V��^�E��e�y�_�u�w�m�F��H����W��_�D��e�d�d�e�g�l�F��s���V��_�D��d�e�e�d�g�l�G��H����V��B��U���w�e�e�d�g�m�G��I����V��_�E��e�e�w�u�w�}�U��I����W��^�D��d�d�e�d�g�m�F��[��ƹF�^�D��d�e�e�e�f�l�F��I����V��_�Y�ߊu�u�e�d�f�m�F��H����V��^�D��d�d�d�d�{�W�W���I����V��_�D��d�e�d�e�f�l�F��I���l�N��E��e�e�e�d�g�m�F��I����W��^�E���u�u�u�w�g�m�F��I����W��_�E��d�e�d�d�g��W���Y����V��^�D��e�e�d�e�f�m�F��H����D�=N��U��d�e�e�e�g�m�F��H����V��^�D��d�y�_�u�w�m�F��I����W��_�D��e�d�d�d�f�m�G��s���V��^�D��e�e�e�e�f�l�G��H����V��B��U���w�e�e�e�g�l�F��I����W��_�E��e�e�w�u�w�}�U��I����V��_�D��d�d�e�d�g�l�F��[��ƹF�^�E��d�d�e�e�f�m�F��I����W��_�Y�ߊu�u�e�e�f�l�F��I����V��_�D��d�e�d�e�{�W�W���I����W��^�E��d�e�d�e�f�l�F��I���l�N��E��d�d�d�d�f�l�G��H����W��_�D���u�u�u�w�g�l�F��H����W��^�E��d�e�e�e�f��W���Y����W��^�E��d�e�e�e�f�m�F��I����D�=N��U��e�d�d�e�f�m�G��H����V��^�E��e�y�_�u�w�m�G��H����W��^�D��e�d�d�e�f�l�G��s���V��_�D��d�d�d�d�f�m�G��H����V��B��U���w�e�d�e�g�l�F��I����V��_�E��d�d�w�u�w�}�U��H����V��_�D��e�e�e�d�g�m�G��[��ƹF�^�E��d�d�d�d�g�l�G��I����V��_�Y�ߊu�u�e�e�g�m�F��I����W��_�D��d�d�d�e�{�W�W���I����V��_�D��d�d�e�e�f�m�F��H���l�N��E��d�e�e�d�g�l�F��H����V��_�E���u�u�u�w�g�l�G��H����W��_�D��d�d�e�e�f��W���Y����W��^�D��d�e�e�d�f�m�F��H����D�=N��U��e�e�e�d�g�m�F��I����V��_�D��e�y�_�u�w�m�G��I����V��^�D��e�d�e�e�g�m�G��s���V��_�D��d�d�d�e�f�m�G��I����W��B��U���w�e�e�d�f�m�G��H����V��_�E��e�e�w�u�w�}�U��I����W��^�E��e�d�e�d�g�m�F��[��ƹF�^�D��d�e�d�d�g�m�F��I����W��^�Y�ߊu�u�e�e�f�m�F��I����V��_�D��e�d�d�e�{�W�W���I����V��^�D��e�d�d�e�f�m�G��H���l�N��E��e�d�d�d�g�m�F��I����W��^�D���u�u�u�w�g�m�G��I����V��_�D��e�d�e�e�f��W���Y����V��_�D��d�e�d�d�f�m�G��H����D�=N��U��e�d�e�e�f�m�G��H����V��_�E��e�y�_�u�w�m�G��I����V��_�E��e�d�d�e�g�m�G��s���V��^�D��d�e�e�d�f�m�G��H����W��B��U���w�e�e�d�f�m�G��I����V��_�E��e�e�w�u�w�}�U��I����V��^�E��d�d�e�e�g�l�F��[��ƹF�^�E��d�e�d�e�g�l�F��I����V��^�Y�ߊu�u�e�e�g�m�G��H����V��^�D��e�e�e�e�{�W�W���I����V��_�E��e�e�e�e�f�m�F��H���l�N��E��d�e�e�e�f�l�G��I����V��^�E���u�u�u�w�g�m�G��H����V��^�D��e�d�d�d�g��W���Y����V��^�D��e�e�d�d�f�m�G��I����D�=N��U��e�e�d�e�g�m�G��H����V��^�D��e�y�_�u�w�m�G��I����V��^�E��e�d�e�d�f�l�G��s���V��^�D��e�e�e�e�g�m�G��I����W��B��U���w�e�e�e�g�m�F��H����W��_�E��d�e�w�u�w�}�U��I����V��_�D��d�e�e�d�f�l�F��[��ƹF�_�D��d�e�e�d�g�m�F��I����V��_�Y�ߊu�u�d�d�f�l�G��H����V��^�E��d�e�e�e�{�W�W���H����W��^�D��e�d�d�e�g�l�G��I���l�N��D��d�e�d�e�f�l�G��H����W��^�E���u�u�u�w�f�l�F��H����V��^�D��d�e�d�e�f��W���Y����W��_�E��d�d�d�e�g�m�F��I����D�=N��U��d�d�e�e�f�l�F��H����V��^�E��e�y�_�u�w�l�F��I����W��^�E��e�e�d�e�g�l�G��s���W��_�E��e�e�d�d�g�l�G��I����W��B��U���w�d�d�d�g�m�F��H����V��^�D��e�e�w�u�w�}�U��H����V��^�D��e�e�e�d�f�l�G��[��ƹF�_�D��e�d�e�d�f�m�F��I����V��_�Y�ߊu�u�d�d�f�l�G��H����W��^�E��d�d�e�e�{�W�W���H����W��^�D��e�e�d�e�g�m�F��H���l�N��D��e�e�e�e�f�l�G��H����V��^�E���u�u�u�w�f�l�G��H����V��^�D��d�e�d�e�g��W���Y����W��_�D��d�d�e�d�g�m�F��I����D�=N��U��d�d�e�d�g�m�F��I����V��_�E��e�y�_�u�w�l�F��I����V��_�E��e�e�d�d�f�m�F��s���W��_�D��d�e�d�e�f�m�G��H����W��B��U���w�d�d�e�f�m�F��H����V��^�D��d�d�w�u�w�}�U��H����W��_�D��e�d�e�e�f�m�G��[���K������0�:�,�9�f�W�W���B���P	��C��U���"�&��0�1�3��������~��[�Oʼ�!�2�'�o�w�}�W��E����V��X��<���-�:��<��>���s���U��N��X��>�:�0�!�8�;�>�������[��V����u�u�n�u�4�3����Y����[��t�����0��'�=�$��6���Y�ƥ�G��EN�U���u�x�i��0�8��������V��E:������!�k�u�w�e�G���Y�����P�����3��1�-�8�	����:����l�N�U���6�;�!�;�w���������r
��T��'���c�!�o�u�]�}�W������U+��X����_�u�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��^�E��d�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�f�l�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�d�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�d�u�}�W���[����W��_�D��e�e�d�d�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��H����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�d�d�f�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��d�w�u�u�w��F��H����W��_�E��d�e�e�e�g�m�F���Y���D��_�D��d�d�d�e�f�l�F��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�E��d�d�e�e�g�m�G��I���F�_�D��d�d�d�e�g�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�d�u�}�W���[����W��_�D��d�d�e�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��H����V��^�E��y�_�u�u�f�l�F��H����V��_�D��e�e�e�e�g�l�[�ԜY���W��_�D��e�e�d�d�g�m�G��I����W�d��U���d�d�d�d�f�l�G��I����V��^�E��d�w�u�u�w��F��H����W��^�D��e�e�e�e�g�m�F���Y���D��_�D��d�e�d�d�g�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�d�y�]�}�W��H����W��^�D��e�d�e�e�g�m�G��H���F�_�D��d�d�d�d�g�m�F��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�d�u�}�W���[����W��_�E��d�d�d�d�g�m�G��I����FǻN��D��d�d�d�d�g�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�l�[�ԜY���W��_�D��d�e�d�d�g�m�G��I����W�d��U���d�d�d�d�f�l�F��I����V��^�E��d�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�F���Y���D��_�D��d�e�d�d�f�l�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��e�e�e�y�]�}�W��H����W��^�D��e�d�e�e�g�m�G��I���F�_�D��d�d�d�e�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�d�u�}�W���[����W��_�E��d�d�e�e�g�m�G��I����FǻN��D��d�d�d�d�g�l�F��I����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�g�l�[�ԜY���W��_�D��e�e�e�d�f�m�G��I����W�d��U���d�d�d�d�f�l�G��I����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�e�e�d�f�l�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��^�E��e�e�e�e�g�m�G��I���F�_�D��d�d�d�e�g�m�F��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��d�d�d�d�u�}�W���[����W��_�E��e�d�e�e�f�l�F��H����FǻN��D��d�d�d�d�g�l�F��H����W��_�D��y�_�u�u�f�l�F��H����W��_�E��d�d�d�d�f�m�[�ԜY���W��_�D��e�d�e�d�f�l�F��H����W�d��U���d�d�d�d�f�l�G��I����W��_�D��e�w�u�u�w��F��H����W��^�E��e�d�d�d�f�l�G���Y���D��_�D��d�e�e�d�g�m�G��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�e�d�y�]�}�W��H����W��^�D��e�e�d�d�f�l�F��H���F�_�D��d�d�d�d�g�m�G��H����W��^�W���u�u�w�d�f�l�F��H����W��^�D��d�d�d�d�u�}�W���[����W��_�D��e�d�e�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��I����W��_�E��y�_�u�u�f�l�F��H����W��_�E��d�d�d�d�g�m�[�ԜY���W��_�D��e�d�d�d�g�l�F��H����W�d��U���d�d�d�d�f�l�F��I����W��_�D��d�w�u�u�w��F��H����W��_�E��e�d�d�d�f�m�F���Y���D��_�D��d�d�d�e�g�m�G��H����V��L����u�e�e�e�g�m�G��I����V��_�D��d�d�e�y�]�}�W��I����V��^�E��d�e�d�d�f�l�F��H���F�^�E��e�e�e�d�g�m�G��H����W��^�W���u�u�w�e�g�m�G��I����W��^�D��d�d�e�d�u�}�W���[����V��^�E��d�e�e�e�f�l�F��I����FǻN��E��e�e�e�e�f�m�F��H����W��_�E��y�_�u�u�g�m�G��I����W��_�E��d�d�d�e�f�l�[�ԜY���V��^�E��d�e�e�e�g�l�F��H����V�d��U���e�e�e�e�g�l�G��I����W��_�D��e�w�u�u�w��G��I����W��^�D��d�d�d�d�f�l�G���Y���D��^�E��e�e�e�d�g�m�F��H����W��L����u�e�e�e�g�m�G��I����V��_�D��e�e�e�y�]�}�W��I����V��_�D��d�e�d�d�f�l�G��H���F�^�E��e�e�d�d�g�m�G��H����W��^�W���u�u�w�e�g�m�G��I����V��_�D��d�d�e�d�u�}�W���[����V��^�E��e�e�d�d�f�l�F��I����FǻN��E��e�e�e�d�g�l�F��H����W��_�D��y�_�u�u�g�m�G��I����W��^�D��d�d�d�e�f�l�[�ԜY���V��^�E��d�e�e�d�f�l�F��H����V�d��U���e�e�e�e�g�l�G��H����W��_�D��d�w�u�u�w��G��I����W��^�E��d�d�d�d�f�m�F���Y���D��^�E��d�d�d�e�g�m�F��H����V��L����u�e�e�e�g�m�F��H����V��_�D��e�e�e�y�]�}�W��I����V��^�E��d�d�d�d�f�l�F��H���F�^�E��e�d�e�d�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����W��^�D��d�e�d�e�u�}�W���[����V��_�D��e�d�e�e�f�l�F��H����FǻN��E��e�e�e�e�g�m�G��I����W��^�E��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�g�m�[�ԜY���V��^�D��d�d�e�e�f�l�F��H����W�d��U���e�e�e�e�f�m�G��I����W��_�E��e�w�u�u�w��G��I����V��_�D��d�d�d�d�g�l�G���Y���D��^�E��d�d�e�d�g�l�F��H����V��L����u�e�e�e�g�m�F��H����W��_�D��d�d�e�y�]�}�W��I����V��^�D��d�e�d�d�f�l�F��H���F�^�E��e�d�d�d�g�l�F��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�e�e�e�u�}�W���[����V��^�E��d�d�e�d�f�l�F��I����FǻN��E��e�e�d�e�f�m�F��H����W��^�E��y�_�u�u�g�m�G��H����W��^�D��d�d�d�d�g�m�[�ԜY���V��^�E��e�d�e�d�g�l�F��H����V�d��U���e�e�e�e�g�l�F��H����W��_�E��e�w�u�u�w��G��I����V��^�D��d�d�d�d�g�m�G���Y���D��^�E��d�d�d�d�f�m�F��H����V��L����u�e�e�e�g�l�F��I����W��_�D��d�e�d�y�]�}�W��I����W��^�E��d�d�d�d�f�l�F��I���F�^�E��e�e�d�d�g�l�F��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�e�e�e�u�}�W���[����V��_�D��e�e�e�d�f�l�F��I����FǻN��E��e�e�d�e�f�l�G��I����W��^�E��y�_�u�u�g�m�G��H����V��_�E��d�d�d�d�g�l�[�ԜY���V��^�D��e�e�e�e�f�l�F��H����W�d��U���e�e�e�e�f�l�F��H����W��_�E��d�w�u�u�w��G��I����V��_�E��d�d�d�d�g�m�F���Y���D��^�E��d�d�d�e�g�m�G��H����V��L����u�e�e�e�g�l�F��I����W��_�D��d�e�d�y�]�}�W��I����W��^�E��d�d�d�d�f�l�F��I���F�^�E��e�d�d�e�f�l�G��H����W��_�W���u�u�w�e�g�m�F��I����V��^�D��d�e�e�d�u�}�W���[����V��^�E��e�d�e�e�f�l�F��I����FǻN��E��e�e�e�e�f�l�G��H����W��^�E��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�g�l�[�ԜY���V��^�E��d�e�e�d�g�l�F��H����W�d��U���e�e�e�d�g�l�G��I����W��_�E��e�w�u�u�w��G��I����W��_�D��e�d�d�d�g�l�F���Y���D��^�E��d�e�e�e�f�l�F��H����V��L����u�e�e�e�g�m�F��I����V��_�D��e�e�d�y�]�}�W��I����V��_�E��e�d�d�d�f�l�G��H���F�^�E��d�e�e�d�g�m�F��H����W��_�W���u�u�w�e�g�m�F��I����W��^�D��d�d�d�e�u�}�W���[����V��^�E��e�e�e�e�f�l�F��H����FǻN��E��e�e�e�d�g�m�G��I����W��_�D��y�_�u�u�g�m�G��I����W��^�D��d�d�d�e�f�l�[�ԜY���V��^�E��e�e�d�d�g�l�F��H����V�d��U���e�e�e�d�g�l�G��I����W��_�D��e�w�u�u�w��G��I����W��^�E��e�d�d�d�f�l�G���Y���D��^�E��d�d�d�e�f�l�F��H����W��L����u�e�e�e�g�m�F��H����W��_�D��d�d�e�y�]�}�W��I����V��_�D��e�e�e�e�g�m�G��H���F�^�E��d�e�d�e�g�l�G��I����V��_�W���u�u�w�e�g�m�F��H����W��_�E��e�e�d�e�u�}�W���[����V��^�D��e�e�d�e�g�m�G��H����FǻN��E��e�e�e�d�g�l�G��I����V��^�E��y�_�u�u�g�m�G��I����W��^�E��e�e�e�d�f�m�[�ԜY���V��^�E��e�e�e�d�f�m�G��I����V�d��U���e�e�e�d�g�m�F��I����V��^�E��e�w�u�u�w��G��I����V��_�E��e�e�e�e�f�m�G���Y���D��^�E��d�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��H����V��^�E��e�e�e�y�]�}�W��I����V��_�D��d�d�e�e�g�m�G��H���F�^�E��d�e�d�e�g�m�F��I����V��_�W���u�u�w�e�g�m�F��I����V��^�E��e�d�d�e�u�}�W���[����V��^�E��d�d�e�e�g�m�G��H����FǻN��E��e�e�d�d�f�l�F��I����V��^�E��y�_�u�u�g�m�G��H����W��^�D��e�e�d�e�g�m�[�ԜY���V��^�D��e�e�d�d�g�m�G��H����V�d��U���e�e�e�e�f�l�F��H����V��^�E��d�w�u�u�w��G��I����W��_�D��e�e�e�e�g�l�G���Y���D��^�E��e�e�d�d�g�l�G��I����W��L����u�e�e�e�g�l�F��H����V��^�E��e�d�e�y�]�}�W��I����W��_�D��d�d�e�e�g�l�G��I���F�^�E��e�e�d�d�f�l�G��I����W��^�W���u�u�w�e�g�m�G��H����V��^�E��e�d�e�d�u�}�W���[����V��^�E��d�d�d�d�g�m�G��H����FǻN��E��e�e�e�d�g�m�F��H����V��^�E��y�_�u�u�g�m�G��I����V��^�D��e�e�e�e�g�m�[�ԜY���V��^�D��d�e�d�d�g�m�G��I����V�d��U���e�e�e�e�g�l�F��H����V��^�E��e�w�u�u�w��G��I����V��_�E��d�e�e�d�g�l�F���Y���D��^�E��e�e�e�d�f�m�F��I����V��L����u�e�e�e�g�m�G��I����W��^�E��e�d�d�y�]�}�W��H����W��_�E��e�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�m�F��I����V��^�W���u�u�w�d�f�l�F��H����W��_�E��d�d�d�e�u�}�W���[����W��^�E��d�d�d�d�g�m�F��I����FǻN��D��d�d�d�e�f�m�G��I����V��^�D��y�_�u�u�f�l�F��I����W��^�D��e�e�d�e�f�m�[�ԜY���W��_�D��e�e�e�e�g�m�G��H����V�d��U���d�d�d�d�g�l�F��I����V��^�E��e�w�u�u�w��F��H����V��_�E��e�e�e�d�g�l�F���Y���D��_�D��e�e�e�e�g�m�F��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�E��d�d�e�e�g�l�G��H���F�_�D��e�e�e�e�f�m�F��I����W��_�W���u�u�w�d�f�l�G��I����W��_�E��d�d�d�d�u�}�W���[����W��_�D��e�e�e�d�g�m�G��I����FǻN��D��d�d�e�e�f�l�F��H����V��^�D��y�_�u�u�f�l�F��I����W��_�E��e�d�e�e�g�m�[�ԜY���W��_�E��e�e�e�d�g�m�G��I����W�d��U���d�d�d�d�f�m�F��I����V��_�E��e�w�u�u�w��F��H����V��_�E��d�e�e�e�g�l�G���Y���D��_�E��e�d�d�d�g�l�F��I����W��L����u�d�d�d�g�m�F��H����V��^�D��e�e�d�y�]�}�W��H����V��^�E��d�e�e�e�f�m�G��H���F�_�D��d�e�d�e�f�l�G��I����V��^�W���u�u�w�d�f�l�F��I����W��_�E��e�d�d�e�u�}�W���[����W��_�E��e�d�e�d�g�m�G��H����FǻN��D��d�e�d�e�g�m�G��I����V��_�E��y�_�u�u�f�l�F��H����V��^�E��e�d�e�d�f�l�[�ԜY���W��^�D��e�e�e�d�f�m�G��I����W�d��U���d�d�d�e�f�m�G��H����V��_�D��d�w�u�u�w��F��H����V��_�D��d�e�e�e�f�l�F���Y���D��_�D��d�d�e�e�g�l�G��I����W��L����u�d�d�d�f�l�G��I����W��^�D��d�d�e�y�]�}�W��H����W��_�E��d�e�e�e�f�m�F��H���F�_�D��d�e�e�d�g�l�G��I����W��^�W���u�u�w�d�f�m�F��H����W��^�E��e�e�e�e�u�}�W���[����V��^�E��d�d�e�e�g�m�G��I����FǻN��D��d�d�e�e�f�m�G��I����V��_�D��y�_�u�u�f�l�F��H����V��^�D��e�d�e�d�f�m�[�ԜY���W��_�E��d�d�e�d�g�m�G��I����W�d��U���d�d�e�e�g�l�F��H����V��_�D��d�w�u�u�w��F��I����V��_�E��d�e�e�e�f�l�G���Y���D��_�D��e�d�e�d�g�m�G��I����V��L����u�d�d�d�f�m�F��H����V��^�D��d�e�d�y�]�}�W��H����W��_�E��d�e�e�e�f�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��_�W���u�u�w�d�f�m�F��H����W��_�E��e�d�e�d�u�}�W���[����V��^�D��d�e�e�d�g�m�G��I����FǻN��D��d�e�e�d�f�m�F��H����V��^�D��y�_�u�u�f�l�F��I����W��^�E��e�d�e�d�f�l�[�ԜY���W��^�E��d�d�e�e�f�m�G��I����W�d��U���d�d�e�d�g�m�G��H����V��_�E��d�w�u�u�w��F��I����V��_�D��e�e�e�e�g�m�F���Y���D��_�E��e�e�e�e�f�l�F��I����W��L����u�d�d�d�g�l�F��I����V��^�E��d�e�e�y�]�}�W��H����W��_�E��d�e�e�e�g�l�G��H���F�_�D��e�d�e�d�g�m�F��I����W��^�W���u�u�w�d�f�m�G��H����W��_�E��d�e�e�d�u�}�W���[����V��^�D��d�e�e�e�g�m�F��H����FǻN��D��d�e�e�d�g�m�F��I����V��^�E��y�_�u�u�f�l�F��I����V��_�E��e�e�e�d�f�l�[�ԜY���W��_�D��d�e�d�d�f�m�G��I����W�d��U���d�d�d�d�f�m�G��H����V��^�E��e�w�u�u�w��F��H����V��_�D��e�e�e�d�g�l�F���Y���D��_�D��d�d�d�e�g�l�F��I����V��L����u�d�d�e�f�l�F��I����V��^�E��d�e�d�y�]�}�W��H����W��^�E��e�e�e�e�g�l�G��I���F�_�D��d�e�d�e�f�l�F��I����W��_�W���u�u�w�d�f�l�F��H����W��_�E��e�e�e�e�u�}�W���[����W��^�D��d�d�d�d�g�m�G��I����FǻN��D��e�d�d�e�g�l�F��I����V��_�E��y�_�u�u�f�l�G��H����V��_�D��e�e�e�d�g�l�[�ԜY���W��_�E��d�e�e�e�g�l�F��H����W�d��U���d�d�d�d�g�m�F��H����W��_�D��e�w�u�u�w��F��H����V��_�E��d�d�d�d�g�l�G���Y���D��_�D��e�e�d�e�g�l�G��H����V��L����u�d�d�e�f�l�G��I����W��_�D��d�e�d�y�]�}�W��H����W��_�D��e�d�d�d�f�m�F��H���F�_�D��d�e�d�e�g�l�F��H����V��^�W���u�u�w�d�f�l�F��I����V��_�D��e�d�e�d�u�}�W���[����W��_�D��d�d�d�e�f�l�G��H����FǻN��D��e�d�d�d�g�l�G��H����W��^�D��y�_�u�u�f�l�F��I����V��^�E��d�d�e�e�f�m�[�ԜY���W��^�E��d�d�e�e�f�l�F��I����V�d��U���d�d�e�e�f�m�F��H����W��^�D��d�w�u�u�w��F��I����W��_�E��e�d�d�d�f�m�F���Y���Z��t�����:�,�9�g�]�}�W��s����c��V	��U����4�!�0��8��������