-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����u
��s�����x�u� �=�%�}����Y����RǶN�����4�u�'�?�4�g�9�����ƴF��C�Bʔ�'�9�g�d�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=C�]���g�d�u�:�.�4��������R
��Y�� ���!�u�:�%�%�)��ԑTӧ��4��_��'���'�0�_�x��)����Y����A��Y��<���'�4�u�;�8�0����s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x��'�8�8�}��Y�Ƙ�Z��E�����u�9�%�3�8�}����Y����k��YחXʓ���!�u�%�}�Ϲ�����V��_�����u�;�7�0�6�9�Z����ƭ�C	�������<�u�4�0�#�<�W�������AF�����߇x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s����R��^��N��� �0�<�0�y�)�(�������R��[����'�'�u�:�<�W�W���Y����6��y�����<�&�&�{�;�f�}�������f(��~#�Uʠ�0� ���y�>��������R
��=d�����u��:��'�4�}�������PF��e�����u�u�!�
�8�4�W��^���9F��X��]���u�4�0�0�{�>����Y����\	��V �U����>�u��w�g��������T��=N��U���u�o�:�!�$�9�������X4��R�����|�_�u�!�%�?��������l��U��Oʷ�:�0�;�_�w�)�����ƨ�A��h�����:�u��u�w�4�����Ƹ�F��R ��1���%�&�n�_�%�5��������G
��QN�����&�u�&�_�w�p����&����G��=N�����9�4�9�o�$�9�������@��V��%���u�!�
�:�>�f�W������l��R ����� �6�<�;�<�8�$���+����e��N�����2�6�u�0�"�3�������Q��Yd��Uʼ�u�0�0��;�z�PϪ��ƾ�G��I�Nʰ�&�u�0� �9�z�P����ƥ�l�R �����!�:�u��#�)�L�������9F�N������4�u�:�2�}����Y����]F��V��ʡ�<�u�&�4�1�4�Z���	Ӈ����=N��Xʷ�u�:�9�1�5�}��������W��NN�����6� �&�:�w�5�W���Y����p*��D�����_�u�0��4�3����Cӏ��U��RN�����!�_�u�u�%�>��������GJ��[��U���7�2�;�u�w�}����+������Yd��U���u�6�u�h�p�z�}���Y�Ʃ�@��E�����1�0��>�w�5����Y�����T+�����u��i�u��}�������F�R ����u�u�0�1�'�2����s�Ʃ�WF��Y�����0��6�;�8�8�L�ԜY�˺�P��A�����3�_�u�x� �}����ӈ��R��X ��%���4�1�4�9�w�4��������VF��CN�����;�!�0�8�3�1�������F��SN�����:�0�u�&�#�8����Y����TF��T�����&�4�{�u�z�+��������]F��EךU���=�:�
�:�6�3����s�ƭ�A�
N��Rʢ�0�u��&�#�<�ϵ�����R
�I�����r�r�_�u��/�K���H�ƻ�V��e��ʴ�1�>�0�0��1�P�������V�=d��Xǣ�:�>�<����W������l��y'������'�>�0�2���ԜY�˺�\	��VN��0ʴ�'�_�u�x�?�2�(���5�ƭ�_ǻC�����
�u�u�9�]�}�Z�������p#��X1�����<�}��|�w�p����������N����>�4��6�]�}�3����Ɗ�p6��N�����'�6�8�%��}�W���0����X��p������&�!�4�~�}�Z����Ʈ�GF��I����u�:�!�8�'�u�W���YӶ��[�V>��Y���u�u�u�u�w�}�ZϷ�Yӕ��l
��^ךU���u��u�k�6�1�[���Y���F�N�U���u�!�
�:�>�W�W���Y���X��[�U���u�u�u�u�w�p�W���Y����_	��Td��U����u�h�u�8������ί�]O�C����&�1�9�2�4�}�W���=���F��N��U���u�u�u�u�w�p����
����\��=N��U���u�u�k�6�~�}�W���Y���F�C�� ���!�
�:�<�]�}�Z�������\<�����9�r�r�2�9�/��ԜY��ƹK�C�����
�u����>�}���T���E��\1��<���u�%�;�u�z�}�Z¨�����%��:��&���:�<�}��$�)�}���T���E��\1��6ʖ�>�u�x�u�z�+����ӥ��g	��C
�����6�;�_�u�z�}�Z�������wF��=N��X���x�=�:�
�w�}�&���T����u��(��0���x�u�u�2�9�/�ϳ�	��ƹK�N��U����h�u�%�9�}�Z����Ʈ�GF��I����x�u�u�:�#�0����Y���F�-��U���
�!��0�>�������K�^ �����9�2�6�u�z�}�W���:���F��\B��U���u�u�u�u�w�}�Z����ƿ�W9��P��U���u�u�u��w�`�W���*����T��T+��Y���u�x�u�;�w�)�(������K�N��1���h�u��u�w�}�W���Y���F�C�����!�
�:�<�]�}�Z���Y�Ɲ�F���N���u�u�u�u�w�}�W���TӉ����h���ߊu�x�u�x�2�9��������t��[�U���_�u�x�0��)�W�������G0��
I�U���0�4�0�u�z�W�W��Y�˺�\	��^N��%����-�u�x�w�p��������}/��X�����x�u�x�=�8��W���Y����G��P�����0�|�u�x�w�p��������%��=N��X���x�=�:�
�w��#�������Z��r ��U���u�x�#�:�<�<�3Ͻ�s���F�A������6�_�u�z�}�1���Y����9F�N��U���0�<�u�4�w�W�W��Y���z(��S����|�u�x�<�w�?���Y���F�N�����u�4�u�_�w�p�W���Y����X��X1�����<�}��&�#�q�W������G��X	�����x�u�u�u�w�}�Iϝ����F�N��U���u�u�x�<�w�.������ƹK�N��U���u�k��
�#��������F�C����&�1�9�2�4�}�Z���Y����F�	N��Y���u�u�u�u�w�}�W���T�ƥ�F��S1�����u�x�u�u�w��W��Y���F�N��U���u�u�u�x�w�(�W���&����Pl�CךU���;�u�0�0�6�8�0�����ƹK��N����;�#�6�;�8�W��������9K�c�����:�<�2�6�:�8�Ϸ�Y�Ư�V��B��&���u�&�&�!�w�8�����ƻ�V��EN���߇x�3�9�u�6�}��������Z��N�����u�:�r�u�%�}�Ϲ�Ӈ��F��^�U���&�!�0�0�z�}����Y����\�C������u�`�m�c�W