-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����0�3�4�6�!�9�Z�������	F��_ �����8�;�x�u�%�:����)����P��g6��*��`�_�x��#�g�E�������V��=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Wǽ�Y����%��N�����4�<�;�9��.��������\��E���߇x��9��0�)�W�������9K�y�����u�;�!� �2�)�W�������/��X�����_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԑT���c��X��Uʁ�<�u�<�0�4�1�����Ƹ�VF��Y��U���0�%�9�!�3�>��������@l�N��U���u�u�:�u�6�5�:���s��ƴF�N��U���>�4��&�6�>�W�������V��_��U���3�<�<�;�$�<�ϫ��Ʈ���Dd�U���u�u�u�u�9�)����YӰ��Z��V��ʧ�;�0�3�:�w�}�ϵ�����P��^ �����u�d�_�x�z�}�W���Y���g���� ���"�9�u�4�4�1��������P	��Q�����u�#�'�u�>�8�Z���Y���F�D<������9�u�&�2�)�Y����ƪ�A��T�����0�!�"�9�w�-����T���F�N�����!�6�:�>�4�>��������@4��C��6���u�&�0�!�y�}������ƴF�N��U���>�#�'�9�4�����Y����P	��Q�����u�<�9�4�'�<�W�������V��T�����u�u�u�u�w�}����
����\��D>�����u�&�;�!�%�:�����ƻ�G��e�����9�6�_�x�w�}�W���Yӭ��CF��_��<���;�=�;�0�w�3����+����A��[�����!�u�2�<�l�p�W���Y���F��EN�����0�<�u��2�>����������B�����=� �1�>�2�}�'�����ƴF�N��U���6�;�!�;�w�2�W����Ư�P
��GחX���u�u�u�u�w�}����4����Z
��V��ʰ�0�,�6�6�2�2�ϱ�Y����C	��G��ʳ�9�0�_�x�w�}�W���YӅ��U ��^���߇x�x�u�u�w�}�W���Ӆ��\��C�����!�6�0�3�4�8�ϻ��Ɓ�pF��DN��ʼ�3�'�0�u�a�?�%���s���F�N��U���&�8�8�'�w�)����Q����A��T�����u�u�|��<�<��������G��q���߇x�u�u�u�w�}��������[	����U���u�=�u�:�1�4����
Ӓ��GF��YN��U���9�0�u�,�8�8�Z���Y���F�D������y�!�0�%�.�W�������\��^�����4�0�4�%�>�9�������F�N��U���0�!�:�u�?�}�6�������V��YN�����>�_�x�x�w�}�W���Y�Ƃ�G�������&�4�>�4�2�4��������u��X�����4�u�0�"�2�}��ԑT���F�N�����<�<�;�&�$�2����Ӄ��[F��^	�������u�=�$�2����	ӏ��]��R
חX���u�u�u�u�#�}�����Ƹ�VF��[����� �0�u�!�>�}��������G�������u�=�!�x�w�}�W���Y�Ƹ�VF��E�����3�6�0�!�#�<�W���
Ӊ��	��C��U���%�;�;�u�$�)���Y���F�N�����6�0�!�!�6�}����ӄ��^��^�����<�=�!�0�8�9�������z��C�����u�u�u�u�w�*��������Z�������<�;�u� �w�.��������Z��C�����0�!�4�1�2�.�Z���Y���F�^ �����0�:�,�}�>�5����Ӓ����R�����4�!�'�6�2�;�����ƿ�_��R
חX���u�u�u�u�5�}�'������9K��C��U���u�u�u�=�w�4��������P��CN�����4�0�u�&�6�9����ӄ��G��R�����u�u�u�u�w�}�����Ʈ�G��QN������{�u�=�w�l��������Z��Y��ʧ�4�u� �_�z�}�W���Y����UF��Z��U���"�9�u�&�#�8�F����ƨ�_��C�����0�!�6�0�1�>����s���F�N��U���u�d�3�4�#�2��������UF��_��<���'�u� �!�'�4�ϼ�Y����S��^חX���u�u�u�u�3�1�Ͽ�Ӓ��]F��S�����=�u�'�2�9�1��������]��XN�����4�0�x�u�w�}�W���Y����_��V�����%�9�!�1�4�8�������KǶN��U���u�u��0�$�>��������P��CN�����4�0�u�&�>�8����Ӓ��G��Q��ʰ�6�%�_�x�w�}�W���YӒ��GF��RN�����&� �0�u�8�1����	Ӓ����Q�����u�;�u�0�#�}���Y���F�N�����0�!�1�7�w�m�Wǻ�����\F��RN�����<�!�'�<�#�/��������R
��@חX���u�u�u�u��8����Ӆ��U ��^��U���6�9�!�:�w�8��������[��S
�����,�4�_�x�w�}�W���YӇ��Z��Y��D��_�x�x�u�w�}�W���Y����^��^��U���u�1�u�&�3�4�W���Y����R��Y�����!�:�u�'�w�2�Ϸ�s���F�N��U���u��a��4�0�������9K�N��U���u��0�%�'�1��������G��B	�����u�:� �0�>�}�W������KǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�9�5�<�Ϸ�����\��=N�����0�0�&�1�;�:���O�ȭ�_]ǻ��U���0�;�8�'�4�.�������F��@��[����%�4�9�]�}��������X��V�����%�4�9�_�w�.�W���ݶ��}��^�����&�{�9�n�w�(�ϩ��Ȝ�T ��T������0�3�6�2�)�Y���B���K��N �����u�'�;�9�#���������JF��[��6����7�_�<�%�/�W���*����F��RN��<���{�6�8�:�2�)�Y���B���F��Y�����!�4�&�4�2�2�}������u��C'�����:�3��9�w�.�WϹ�����l�N�����9�6��6�8�}�W�������V��V ��U���:�f�o�u�l�}�Wϵ�����G��RN����2�'�n�u�'�/�_���Yӵ��C
��[��U���&�1�9�2�4�W�W���+����A��[��U���7�:�0�;�]�}�W�������\��YN�����0�}�m�1� �)�W���Y���fT��d��Uʦ�:�3��!�m�2�ϭ�����V��X����|�u�x�u�e�s�}���Y����G/��R������9�n�_�%�5��������g*��QN�����;�0�%�:�1�����
���K��R��ʡ�0�%�%�9�9�}����Y����Z��_�����4�!�;�0�'�0����
Ӓ����VךU���<�u�=�&�1�1�Yϊ��Ʃ�@��DN�����3�9�&�>�8�}����ӂ��R��C�����x�1�!�u�6�5�W�������C��R�����<�<�;�u�9�}��������^��d��U���!�%�u�:�1�����	����R��Y	��ʼ�u�;�0�0�w�<����Y����G	�d��X���0�<�,�>�8�;�4���)����V
�������4�2�u�0�>�8�W���:����p��g��1���,�4�2�
�y�}�Z�������A��C�� ���:�9�u� �'�/�ϭ��ƾ�]��=N�����4�!�>�0�>�$����:����Z��R��U���3��9��'���������Gl�N��U���u�u�u�u�w�}�W���Y���F�S��6���3�4�6�<�2�8���s�ƿ�T�������0�:�,�o��+�A���&����U��X����_�u�u�u�w�}�W���Y���F��-�����3��4��%�$����0����]�������:�>�4�!�%�f�}���������D�����6�<�0�o�5�2����C�ƪ�_��=N�����9�&�0�1�3�/����Y����T��F����!�u�|�h��)����D���O��C� ��d�_�u�&�0�<�W�������R)��T�����:�<�
�0�#�/�D�������V�S�����'�u�k�r�p�f�Wϭ�����@4��S*������%�u�u�#�����&����\�N�����u�|�o�u�8�5����G����]ǻ�����&�:�3�<�>�3�W�������T��S�����|�o�u�:�?�/�W���^���K�d\�D���x�u�=�u�%�9�����ƥ�@����U���a�u�9�8�9�}����Y����V��C�����3�u�x�u�c�s�[ϩ�����R�N�����:�4�u�<�$�}�4�������]��R��U���;�,�:�0�:�/�}���TӀ��P��Y�����u�:�3�!�>�)�W���Ӕ��A��Y�����7�3�'�u�2�>�Ͽ�Ӓ��^Hǻ�����!�>�:�3��4�������R
�
N�N���&�2�4�u��8��������@��R
��Aʱ�"�!�u�|�m�}�������A��U��Xʆ�`�x�_�u�$�:����?����c��R'�����u�u�;�<�9�9�E�������V�S�����'�u�k�r�p�f�Z���K����F��P ��U���4�!�=�&�����Cӓ��Z��SF�U���;�:�e�u�j�u����
���V�N�U��{�_�u�<�9�1��������@��g��G�� �&�2�0��m��������\������h�u�e�|�w�p�"��I����Z��[N������4�0�;�>�8�W�������V�N�����u�|�o�u�8�5����G����]�N��D��_�u�<�;�;�.����=����c��N����0�}�a�1� �)�W���C����G��DN��U��|�u�x��b�p�}���
����_F��X�����;��%�e�m�.����Q����\��XN�U��}�!�0�&�j�}�G���Y����W�=N�����9�&�:�3�>�4����	�����Y��G���:�;�:�e�w�`�_������F�G�X���g�{�_�u�$�:����:����p��T�����1�&�:�3��)��������N��_��U��r�r�n�x�w�o�Y�ԜY����R
��t�����6�<�0�o�$�:����:����|��E�����h�}�!�0�$�`�W��P���5��_װU���u�;� �0�#�<�W���Y����_�������4�!�'�!�2��'ϼ�����]��R��ʴ�0�;�!�u�z�}��������Z��=��Fئ�u�4�!�<�"�8����Y�ƿ�A��d�����<� �0�>�2�}�ϭ�����F��D�����&�w�'�0�l�}����������GN��U���0�3�6�0�#�4���
����_F��L�� ���_�u�!�'�5�)�W���	Ӊ��@%��Q�����<�0�o�&�0�<�W���[����]ǑN����>�&�2�!�%�W�W�������@��Y
װ���;�u�x�u�%�<�Ͽ�����V��e�����4�6�_�u�w�/����Q����_��\GךU���0�<�_�u�w�}�Ϭ�
����V��=�����9�|�!�0�]�}�W���Y����G��t��%���u�h�&�0�#�/�4���B���F��Y
���ߊu�u�;�u�%�>���s���%��V�����4�1�0�&�1�/����;����Q��SN��U���0�4�<�;�8�3�W���Y����@��=N�����&�}�4�%�2�1�^�������9F������;�
�1�0��0�����Ƹ�VǻN��U����0�!�u�?�}����
�ƪ�AF��RN�����6�0�3�6�2�)����T����JF��S��U��u�:�!�0�w�}�W��Y����T��U��U���&�=�&��]�}�W���Ӎ��V��X�����'�h�f�u�9�}�%�������_��_��U���u�u�&�0�3�9����Y����V��RF������}�m�1� �)�W��U���F�D��7����9�0��#�/�1�������9F�N��Xʖ�0�!�u�=�w�9����Y����G��D�����:�3�<�<�9�}�����Ʈ���^ ��D��!�u�=�_�w�}�W������V��^������4�0�;�w�}�Wϻ�
���X)��E�����6�:�u�u�w�3�W���
����p��N��U¾�#�'�9�6��>����Y�ƭ�WF��R�����9��%�|�#�8�}���Y���@4��S/�����u�h�'�&�-�u�'������F��@ ��U��y�e�u�u��.�1�������V��V���ߠu�u�u�x�w�/��������W��D�����=�u�<�&�w�2��������_	�������&�;�u�=�w�3����s���F���ʺ�u��4�0�9�}�W�������F�N�����1�1�'�&�w�`�����ο�[��~ ��Mʱ�"�!�u�d�{�m�L���Y����]��QUךU���;�u�3�_�w�3�W�������9l�C�����u�=�u�:�1�4����Y����A��e/��]��>�|�_�u�z������Ư�V ��T��ʴ�1�1�9�4�1�2�W���Y����Aǻ�����}�4�%�0�;�t�Wϼ���ƹF��QN�����
�1�0��:�1�4���Y����9F�N��'����!��!�k�}�4�������A��X1�����'�&�0�1�3�/����B���F��e��1����!�<�0�k�}�%���=����F��N�����<�n�u�0�3�-����
��ƹK�t�����0�!�<�u�'�8�W������"��C��ʻ�-�u�:�3�>�4����
ӊ��V�N���ߊu��0�3�4�8���
����WN��R����� ��%�}�b�9� ���Y���l�D-�����9�4�i�u�>�3�ǭ�����G��C>����u�:�;�:�g�t�}���	����@��V�����|�u�7�2�9�}�WϷ�Y����]��S	��&���9��>�u�?�3�W���Y���c��[��U���u�'�6�<�9�1����Y����c��R'�����=�!�<�u�>�8�W�������G��T�����;�<�2�u�w�}�Z�������9F�N��3���!�=�&���-�G��Y����@��\����!�u�|�_�w�}�W�������R��Y>�����h�&�'�6��<��������9F�N��3���!�=�&���-�E��Y����P��V�����0�n�u�u�w�.����)����z��G�I����4�!�=�$��'���K���F�C�����%�%�9�;�w�)��������VF��E�����<�<�2�7�#�8�Ϫ�Ӥ��~F��SN��ʑ��m�u�9�4�W�W���Y����U ��[�����u�h�&�:�1�����s���F�>�����0�:�<�<�6�}��������GF��XN�����!�0�1�9�6�9����Y�����R�����!�<�0�u�j�.��������G]ǻN��U���0�3�6�0�#�4����D�ƿ�\��^�����%�e�_�u�w�3�W���s�Ʃ�WF��X���ߠ_�u�u�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǻC�!����9�<�9��9���<ӄ��P��Y�����!�&�4���e�[Ͻ�����A��Q��ʸ�9�<�9�_�w�p�W���Y����U��C��[���x�u�!�<�w�2��������Z��a�����y��'�0�w�}��������Q��g)��[���x�u�u�u��2�W�ԜY���W��qN��U�ߊu�x�u�d��}�ϝ�Y���F��e��U���u�u�u�0�]�}�Z���4���rL��N�U���u�h���w�p�}���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�Uʘ�9�<�9��3�.�Cכ�Y����XF��=N��U���%�;�;�u�$�i����Y����V��^��U���u�u�����W���Y���F��^ �����o�u�n�u�w�}�Wϟ�,����a#��N��U���o�<�!�2�%�g�W��Y���F��e+��U���u�u�u�u�w�g�������F��=N��U���u� �����6���+����g#��N��U���o�7�:�0�9�g�W���*��ƹF�N�� �����
����(���<����c2��aN����;�u�h�w���U�ԜY���F��~ ��!���u�u�u�u�w�}�������"��r-��N���u�u�u����2���Y���F�N�����'�o�u�n�w�}�W���;����F�N��U���u�o�<�!�0�/�M���B���F�,��;���u�u�u�u�w�}�Mϭ�����	[�s'��6���_�u�u�u�w��%���+���F�N��U���0�0�u�h�f�W�W���Y�Ə�a4��y=��'���u�u�u�u�9�8����D����F�N��6���u�u�u�u�w�}�W���Y����T��S��N���u�u�u���}�W���Y���F�N�����6�:�u�h��n�1���?����uD��N��U�����u�u�w�}�W���Y����Z��P��O���n�u�u�u�w��;���+����a#��N��Oʼ�!�2�'�o�w�f�W���Y����c+��r<��U���u�u�u�o�>�)����C����9F�N��U�����u�u�w�}�W���Cӄ��l��C��O���w�e�e�e�g�m�G��Y���F��e+��U���u�u�u�u�w�g�������F��=N��U���u��
���}�W���Y�����^ ��O�����w�_�w�}�W���<����g2��yN��U���u�u�!�<�0�g�W͎�-����]ǻN��U����
�����:���Y����G��PN�UȆ����w�]�}�W���Y����~)��N��U���u�u�u�!�>�:�M���*����l�N��Uʀ����u�w�}�W���Y�ƿ�A��T��W�����n�u�w�}�Wϋ�<����g#��h*��0���o�&�'�;�w�`�U���)����gD��N��U��� ����w�}�W���Y����@��Y	��H����a�w�n�w�}�WϮ���ƹF�N��9���u�u�u�u�w�g����
����_	��TUךU���u�u�u�u�w�}�W���Y����]F��C
�����
�0�!�'�e�}�������9F�N��U����u�u�u�w�}�MϷ�Yӕ��l
��^�����'�g�u�:�9�2�G��Y���F��t!��U���u�u�u�o�8�)��������l��C��G���:�;�:�e�l�}�W���YӤ�F�N��U���o�<�u�&�3�1��������AN��
�����e�n�u�u�w�}�5���Y���F�N����&�1�9�2�4�+����Q����\��XN�N���u�u�u���	�W���Y���	F��CN�����2�6�#�6�8�u�@Ϻ�����O��N��U����u�u�u�w�}�W���Y���@��[�����6�:�}�b�3�*����P���F�N��U���u�u�u�u�w�}��������T��A�����b�1�"�!�w�t�}���Y���c%��N��U���u�u�u�;�w�)�(�������P��Z����!�u�|�_�w�}�W���:����F�N��U��� �u�!�
�8�4�(������F��@ ��U���_�u�u�u�w��%���Y���F���U���
�9�2�6�]�}�W���Y����j)��N��U���u� �u�!��2��������U��X����n�u�u�u�w��%���8����F�N��Uʦ�1� �:�<�l�}�W���Yӥ��a?��d-��!���o�:�!�&�3�(����B���F�!��:���u�u�u�u�m�4�Wϭ�����Z��R����1�"�!�u�~�W�W���Y�ƍ�f+��rN��U���u�u�;�u�#�����&����\�
�����e�n�u�u�w�}�4��� ����F�N����&�1�9�2�4�+����Q�ƨ�D��^����u�u�u� ���9���Y�����D�� ���<�n�u�u�w�}�:���*����f2�N����&�1� �:�>�f�W���Y����e#��{!��U���u�o�:�!�$�9������ƹF�N��;�����u�u�w�g����
����_	��TUךU���u�u�����2���-����F��C
�����6�_�u�u�w�}�6���+����v%��T�� ���!�
�9�2�4�W�W���Y�Ə�rW�N��U���u�u�;�u�#��������F�N��4���u�u�u�u�w�}��������\��d��U���u��� ���W���Y�ƥ�F��S1�����n�u�u�u�w��5���Y���F�N��Uʦ�1� �:�<�l�}�W���Yӥ��F�N��U���o�<�u�&�3�(����B���F�-��U���u�u�u�u�m�4�Wϭ�����T��=N��U���u�����}�W���Cӏ����h�����_�u�u�u�w��#���Y���F���U���
�9�2�6�]�}�W���Y����F�N��U���u�;�u�!��1����s���F�t+��9������u�w�3�W���&����Z��N��U�����u�u�w�}�W���Y���@��B����u�u�u�u��	�W���Y���F��^ ����� �:�<�n�w�}�W���+����%��e7��U��<�u�&�1�"�2���Y���F��d:�� ����u�u�o�>�}��������P]ǻN��U�����u�u�w�}�W������G��[���ߊu�u�u�u���W���Y���\��YN�����9�2�6�_�w�}�W���*����F�N��U���;�u�!�
�;�:��ԜY���F��c#��U���u�u�u�u�9�}��������l�N��Uʇ��u�u�u�w�}�W����ƿ�W9��X	��\�ߊu�u�;�u�8�-����B���F��P ��U���9�u�u�!��2��������T��S�����|�_�u�u�>�3�ϭ�*�����h�����0�!�'�d�w�2����I��ƹF��^	��ʦ��#�o�&�3�1��������AN��
�����e�n�u�u�$�:����)����	F��S1�����#�6�:�}�`�9� ���Y���9l�U���ߊu�u�x��w�5�W���M˃�rF��SN�����u�;�u�<�2�4�ϭ�����V ��RN��ʘ�8�9�<�9�2�s�W���T�Ƙ�VF��D��U����=�&�:�2�-�����ƿ�R��U�����=�u�u�1�2�s�W���T�Ƙ�VF��E�����&�'�2�&�2�8�W�������[��^ ��U���%�!�_�u�w�p�W�������c��R'�����u�;�u��2�;����)������Z�����0�u�;� �$�W�W���8����[��C
�����
�0�!�'�%�.����?����c��R'�����y�e�|�u�z��G��Y����q5��R�����9�2�6�#�4�2�_�������p	��Q*�����%�e�d�|�l�p�W��W��ƓF�C�����;�&�:�3�>�4����	���F����U���0�u�;� �y�}�Wϭ�*���F��S1�����#�6�:�}�2�4�ǭ�����P��C>�����&��#�9�9�)�W���:����`��CG��Sʯ�'�&�>�:�1�����B���`R�� dךU���&�a�0�-�m�9����s���T��E�����_�u�u�u�4�.����D����9F�N�����1�'�2�h�w�q�W���YӇ��TF�_�U���u�4�!�'�$�)��������V��CN��U���&�y�u�u�w�<����
����R��E �����!�:�!�;�w�c�U���:����F�N�����!�h�u����U�ԜY���Q��T��U��d�_�u�u�w�/���Y��ƹF������u�k�w���	�[���Y����R��^ ����u�y�u�u�w�>��������V�	N����u�u�'�2�j�}�[���Y����R��
P��Wٓ������q�W���YӋ��TF�_�U���u�8�9�6�%�$����Y���l�N�����1�'�2�h�w�q�W���YӖ��G��S���e�e�e�e�g��}���Y�Ƽ�V�	N����u�u�0�
�8�3��������X�d+��8���w�_�u�u�w�8�(������+��|L�U���u�&�9�%�#�8���YѶ��g#��BךU���u�&�
� �#�`�W͓�5����l�N�� ���%�!�0�;�3�)����G�Ă�l6��s+��Y���u�u� �0�$�0�W���[����D�N�����u�4�}�u�w�}����D�Ɵ�^��t�����u�u�u�k�$���ԜY���QF������u�u�u�6�j�}�4���U���F��V�����k�r�r�_�w�}�W������	��R��H���e�|�_�u�w�}����D����G��DN��U��|�_�u�u�w�>���Yۉ��V��
P��E���_�u�u�u�6�/�������A��d��U���8�9�&�2�>�}�I���^���F�V����u�%�;�_�w�}�W������	��YBךU���u�4�'�6�$�2���Y����l�N�����&�2�:�!�j�}����s���F��
P��%���y�u�u�u�'�)��������GF����ߊu�u�u�4�#�/�������	��YBךU���u�#�'�9� �`�W������F�B �����"�h�u�%�9�W�W���Y����J	��S����y�u�u�u�'�2���Y����l�N�����1�u�k�w�f�m�G���s���F��B����u�e�e�w�]�}�W�������]��S�W��w�_�u�u�w�8�F��Y���9F�N����h�u�d�y�w�}�WϽ�����W�	N��R�ߊu�u�u�0�f�`�W��U���F��R�H���d�y�u�u�w�>���Y���9F�N�����'�<�u�k�p�z�}���Y�Ư�^F�I�Y���u�u�6�6�%�}�I���^���F�T��H���d�y�u�u�w�>��������Z�	N��R�ߊu�u�u�&�6�`�W��U���F��D�� ���0�h�u�e�{�}�W�������X�I�U���u�'�!�u�i�z�P�ԜY���A��[�����;�h�u�e�{�}�W�������X�I�U���u�'�!�!�;�`�W��U���F��D��H���e�|�_�u�w�p�W�������[��d>�0ʺ�!� �_�u�w��������F��P ��]���9�}��0�1�(�P�������p	��Q=�����:�;�:�>�8�;�$�������F��SN������9�<�9��9���<��ƹK�g�����u�=�u� �'�)��������G��N�����%�%�9�;�w�)����
ӎ��VF���� ���'� �<�2�w�p�W����Ʈ�G��YN������a��7�8�6��������r%��d>�0ʷ�:�>�u�%�8�8�Ǎ�����_�N�����u�u�<�u�>�4�����Ο�^��t��U���;�u�u�u�$�2��������VF������4�6�_�u�w�3�W���s�Ʃ�WF��X���ߊu��0�3�"�}�Jϭ�����R
��^����1���_