-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B ��X��ģ�1�x�u� �?�/�W���Y����Al�!�����9��:�0�#�}�/���L����9K�s��O���;�u�e�d�p�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d�U¶�u�e�f��'�/����7����]��~ �����;�&��'�8�<����T�ƍ�_F��P��U���0�#�1�x�w�<����ӯ��G��R ��U���0�;�9��1�/�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�x�u� �'�.�M��Y�Ƙ�Z��X�����u�&�&�8�;�}�W���&����PF��N�����u�4�u�4�8�)��������GHǶN��!���u�4�u�0�"�8�W����ƅ�z(��YN��U����!�u�0�w�}�1ϩ��ƭ�X����U���:�!�x�u�w�2�������2����U���:�!�<�u�2�}�Ϫ�Ӆ��_��=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W��������V��=N�����0�0�&�1�;�:���O�ȭ�_]ǑR �����$�4�:�!�1�4�W�������PNǻ�����:�!�u�u�#�4���Y���]��X�����4�%�0�9�w�}�W���Y����Z��C
�����n�u�&�4�6�3�W���Y���F������9�2�6�_�w��������F�N��Oʺ�!�&�1�9�0�>�^����Ɖ�u��B��N�ߠ4�6�<�0�#�/�W���Y����B ��X��ʼ�_�u�&�2�6�}�3���6����_F��D�����6�o�u�e�l�W�W��2����\��_��3���4�!�<� �2�6����Y����]��N����� �0�>�0�w�;��������P
�N�����u�&�w�'�2�f�}�������F��Z����� �o�&�'�9�f�WϿ�����G��V�����!�:�u��#�����Y�ƿ�T��������;� �n�]�8��Զs�Ɗ�Z��X�Uʥ�:�0�&��:�1�4���s�Ʈ�T��N�����<�<�2�0�0�u����������Yd��U���&�4�4� ��1�K���=����]]ǻN�����3�_�u�;�w�/����Y����u
��dךU���!��!�i�w���������9l��Y
��!��