-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����;�!�:�!�8�s��ԑTӧ��[	��$��ʔ�8�'�4�_�z������Ɯ�\��CT��-���`�a��x�w�<����Oӫ��T��d����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z���P����F��G������!�:�4�w�3��������p	��X�����x�u�9�u�>�5�ό�
����Wl� �����9��&�'�:�3�ϗ�����_F��Q�����;�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���6��G��O���=�&�3�9�w�0��������[��X �����;�!�3�'�#�8��������_F��T�����x�u�u�u�w�}�W�������]��Y��Uʐ�6�u�'�6�$�4�ϫ��ƻ�_
��V�����:�;�6�;�%�1�Z���Y���F�U������0�6�;�%�1����Ӓ��_��_�����:�u�=�u�%�>����ӓ��GF��R חX���u�u�u�u�6�>����������S��ʷ�u�!�'�y�?�*����Y����V��_�����9�!�:�_�z�}�W���Y����Z
��T�����y�4�1�"�6�}��������GF��V��U���u�&�1�3�%�)���Y���F�N�����4�<�;�u��}��������_��DN��ʦ�4�!�%�4�2�;�Ϫ�ӈ��Gl�N��U���u�u�:�!�8�}��������V
�������u�:�&�4�#�4�ϰ��Ư�_��V���߇x�x�u�u�w�}�W���
�ƿ�V��E��ʳ�'�0�!�0�4�3��������G	��P ��ʡ�0�6�'�0�#�p�W���Y���F��[�����;�4�1�%�2�<�ϸ�Ӈ��V��Y�X�߇x�u�u�u�w�}����
����A��Y�����u�=�u�:�#�2�W����Ƥ�DF��T��ʼ�6�0�0�!�#�8�Z���Y���F�T�����3�'�0�6�w�8�W�������Z	��=C�X���u�u�u�u�w�� ���:����z��O(��!�����u�&�$�?�����ƪ�\��_�� ���;�u�=�&�]�p�W���Y�����X�����2�&�;�u�?�}����=����V ��V��Uʁ�<�u�&�1�9�}�Ϫ��Ƹ�Vl�N��U���u�u�:�3�>�4��������CF����U���'�u�!�4�3�8�Ϥ��ƣ��������_�x�x�u�w�}�W���Y����[��t�����0��'�=�$��W����Ƹ�VF��Y��ʠ�<�u�3�!�2�>�������F�N��Uʶ�0�3�6�0�#�.����Y����V��T�����=�&���8�}�����Ƹ�VF��O�X�߇x�u�u�u�w�}��������V��Y�����0�9�u�=�$�?��������R��T�����!�&�:�9�w�-��ԑT���F�N�����9�!�;�u�2�2�Ϸ�Y����@F��RN�����!�u�=�u�2�)�:���Yӯ��G��=C�U���u�u�u���5�ϸ�����WF��[N��U���u�:�3�<�>�3��������VF��RN�����!�x�u�u�w�}�W�������Z��E�����=�;�&�<�?�.�4�������K ��c��8���u�=�;�!�>�}�6�ԑT���F�N�����&�4�9� �#�1����Y����[��T�����1�4�9�:�w�)�W�������Z	��C��U���u�u�u�,�;�.�}��T���F�N��!���%�%�9�;�w�8��������`��C>�����9�1�!�u��%�:�������F��[��X���u�u�u�u�w�.����Ӓ��@%��T-�����<� ��0�|�l�}��T���F�N��!���%�%�9�;�w�8��������`��C>�����9�1�!�u��.��������]ǶN��U���u�u�&�4�4�5��������WF��]�����u�,�9�&�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=d�����,�<�0�y� �/�L�������V��D�����6�d�c�{�;�f�Wϫ�ӏ��VH��Z�����1�4�9�_�w�.�W���݈��V��h��[���n�u� �0� �/�Y���7����_��R��Ĵ�9�_�u�&�w�2��������G��V�����!�'�4�9�]�8����Y����G"��g�� ����;�'�9�>�W�W������F��Z��6���o�<�u�!��2���s���@4��C��U���o�<�u�:�;�<�L�ԜY�ƿ�[��~ �����!�o�<�u�9�4��������[��u��X���:�;�:�e�l�}�Z��W��ƹF��{�����0�3�;�0��/����8����Z��Y�����d�u�:�;�8�m�L���T����TǻN��=���0�!�:�3��9����-����r%��� ���2�0�}�d�3�*����P���3��_�U���&�4�6�,�;�.����6�����B �����}�u�:�;�8�m�L���T���9l�N������4�0�4�>�}�W�������R��N�����'��4�0�m�4�W���������Z>�����!�x�u�:�9�2�G��Y�˙� H��=d��Uʦ�0�!�4��6�8�������	�������n�u�u�&�2�)��������GF��X�� ���2�0�}��:�5��������W	��C��\���x� �f�d�]�}�Wϭ�����G%��TN����7�:�0�;�]�}�W�������@��C8�����u� �u�:�;�<�L���Yӕ��_��V�� ���u� �u�;�>�3�ǵ�����P6��D�����u�:�;�:�g�t�W��,���l��SN�����0��:� �>���������A��C�� �����:�u�%�>�3�������Z��Y��ʼ�_�u�x�u�8�/�����ƣ��������<�;�9�4�2�>����Ӓ��A��T�����4�x� �u�9�)�������F��P ��U���9�u�u�:�;�<�!�������W	��C��\��u�:�=�'�w�c����P��ƹ��Y�����!�'��%�w�}����������RUװU���u�=�u�,�;�}�����ƿ�R����G���=�&�4�9� �}�Ϫ�Y����_�������8�9�!�_�w�p��������GF��S�����'�u�=�u�2�)��������@��[�����:�&�4�!�<�<��������F��Y��Oʠ�&�2�0�}�w�2����I����D��^�D���u�x�m�m��1���K���@��V��6����6�0��"�)�Mϫ�
����WN��S�����|�o�u��;�����:����z��N��X��m�u�&�2�6�}�'�������^F��B �����}��8�=�$����Y����G	�N�Uº�=�'�u�k�p�z�L���T����TǑN�����u��-��4�5���������^	��¾� ��4�0�>�.�FϺ�����O�
N�����&�h�u�e�~�}�Z�J����F��P ��U���-��6�=�$�����Cӄ��_��T�����n�u�&�2�6�}�9���4����R��B��%���u�u�:�9�6�}�JϪ���ƹ��Y�����!�4��4�2�(�;���Cӓ��Z��SF�� ���4�0�<�&�f�9� ���Y���F��C����u�e�|�u�z��D��s���@��V��6����4�0� ��1����	����\	��V ��Hʳ�9�0�_�u�>�3�ϭ�����G%��T:����7�:�0�;�m�}����B����Z��[N�����4��4�0�"���������Q	��R��O���4�&�n�u�$�:����+����A��[����7�:�0�;�m�}����B����Z��[N�����=�&��!�6�4�;���Cӄ��_��T�����0�_�u�<�9�1��������V)��{��Oʠ�&�2�0�}��0��������Z��N�����u�|�o�u�8�5����G����]�C��F��_�u�&�2�6�}�%�������_��[>����7�:�0�;�m�}����B����Z��[N�����=�&��!�6�4�;��������[��U��3�9�0�_�w�4����
����c��R!��9����0�o� �$�:����7����_��V�����d�1�"�!�w�t�M�������@F�I�\���x� �f�d�]�}�����ƿ�R
��N����� ��0�<�2�g��������F��@ ��U���o�u�:�=�%�}�I���^���3��d�����4�u��9��0����Y�Ʈ�\
��YN�U���&�n�_�u�#�/����Y����\��C���ߊu�x��&�%�}����������Y�����:�u�0�2�3�*�������� ��ZN������'� �<�$�.�W���Ӓ��9F�N�� ���2�1�9�,�>�}����s�ƭ�G��B�����u�3�&�0�#�/�'���Cӕ��]��^�����w�_�u�x�w�<�ϭ��Ƹ�R��_�����<� �9�&�3�8��������A��X�����<�0�u�;�8�2�ϭ�����9F�N�����<�9�=�9�w�4�ϸ�މ����^ �����0�{�u�4�#�4��������\ ��~
��Oʦ�2�4�u�&�u�/���YӇ��A��C�����:�u��9��>��������V6��RT�����9�<�u�!�"��}���T�Ɯ�V��CN�����=�&��!�6�4�;�������A	��U��ʸ�'�0�u�<�?�)�Ϯ�	����VF��P �����x�u� �&�3�}��������JF��EN�����u� �%�&�$�W�W�������VF��R��ʦ�4�6�=�&��)����5����C��D�����&�w�'�0�l�W�W�������@��C�����x�=�:�
�>�8��������9F��E�����4�%�0�9�~�}���������E�����1�0��8�;�������ƹF�C�%���9�;�u��$�<�Ϫ�Y����A	��^ �����u�u��&�6�)����E�ƿ�V��E�U���u�<�u�&�2�)����	�Ƹ�VǻN��U����9�u�h��)����D�Ƹ�F�=N��U���;�u�3�_�w�}�W�������_��^ ��:���<�0�i�u��1�4�������F��RUךU���u��9��:�1����Dӕ��_��T��6���!�h�&�4�4�$��������]��G�U���u�x�u�0�6�1�W�������]��N��Uʦ�0�!�4��6�8��������_F�����u�u�u�&�2�)��������CF�����u�u�u�&�6�>����6����_��R��I���4�&�n�_�w�}�W��:����_����U���9�4�u�:�#�2�W�������F��PN�����e�_�u�u�w�;���������Yd��U���u�x�u�:� �}����Ӑ��Z��C��U���&�j�u�3�$�q����Ӈ��R
��[�����u�u�u�u�z�}�ϭ�����G6��RN��U���0�!�1�<�9�/�W���Y����A��V�����{�u�u�u�w�4�_�������R��V��U���u�:�u��$�<�����Ƹ�VǻN��U���u��&�4�#�<����	���G��d��U���u�u�&�4�4�5��������W2��GN�U���0�_�u�u�w�}�W������N��_��U��3�9�0�n�w�}�W�������U]ǻN��U����u�'�u�9�)�Ϯ�����Z��D�����u�u�0�&�]�}�W���Y����P6��D�����<��8�u�j�)���Y���F�N��ʢ�u�:�0�"�#�}��������R��YN�����_�u�u�u�w�;��������_��N���ߊu�u�u�u�w�����D�Σ�[��S����|�_�u�u�w�}�W�������c��R!��#���1�6�u�h�#�(�L���Y����������u�u�;�u�1�W�W���Y���p��B��ʦ�4�6�,�9�$�2����
����@/��RF����u�u�3�&�3�8�F�������F�N�����6�,�9�&�8�3�W������p��R�� ���;�!�_�u�w�}����Y���F��t��6���0�� �!�k�}�4���:����@%��Y��U��u�u�u�0�3�4�L�ԜY���K��V�����u��4�0�4�(�W����ƿ�W
��GךU���u�3�&�1�2�o�^Ϫ����F�N������6�8�i�w���������9F�N�����u�u�u�u�$�5�������F��_��4���8�~�&�=�$���������F�N��ʼ�n�_�u�u�w�p�4���������O�����&��6�8�"�4�ϭ����l�N��X���:�<�0�!�6�}�Ϸ�����Z��D ������4�0�6�"�}�ϭ�����[��E��G���&�=�&��4�8����W����[��N��U���u�&�1�;�w�8����Y����Z��^ �����!�4��4�2�>�����ơ�A��^�����'�u�!�<�w�8�Ϫ�Y����]��#��[���u�u�x�u��%�:�������P�������,�u�6� �;�$����������V
��ʢ�0�0�<�u�?�(�ϼ�Y����P��Z�����=�&�u�u�w�p�W����Ƽ�C��Y�����{�u�u�u�>�u�>���Q���G��=N��U���u��-��4�5�������F��C��%���0�~�}��6�8��������@6��D�����0�!�=�2�z�}�������F�G�U���u�0�&�_�w�}�W���7����R��V�����u�h�&�0�#�<�'�������^F�D>�����6�0�0�!�]�}�W����ƥ�lǻN��U����!�'�<�2�*�����Ƣ�K��v-��U���&�u� �u�?�(�ϼ�Y����G��N�����&�0�!�4��<����<�ƥ���^�����_�u�u�u�z�.��������@��C"��U���9�&�:�u�'�<��������Z��DN�����'�!�4�u��:��������]��q������{�u�u�w�.��������@��C+��I����-��6�?�.�6���ۍ��^6��D�����u�:�;�:�<�(�'���������P�����3��1�-�8�	����:Ԋ��T��R�����=�&��0�1�3��������~'��=d��U���x�u�'�4�2�)�ϸ�����}��z������!�6�_�w�}�W���
����~��_��:���;�u�=�;�w�}�W���
����~��_��:���6�u�h�&�2�)��������P��=N��U���;�u�3�_�w�}�W��Y����_�������6�=�&��#�3��������G��=N��U����-��6�?�.�8�������Z�D ������4�0� ��f�}���Y���6��R��ʇ�&�4�!�4�4�<�ϝ�����@��C8�����2�<�u�:�4�0�����ƪ�AF��RN�����%�%�9�;�w�)����ӥ��P6��D��ʷ�9�"�_�u�w�}�Zϝ�����@��C8�����=� �1�4�$�/�W���Y����F��D�����6�6�u�&�2�)�Y���ӕ��F
��V��U���0�!�4�,�#�0�W�������@��C8�����8�_�u�u�w�p��������]��RN�����:�0�6�0�1�>����Y����R
��[��U���=�!�<�u�8�)�������p��g��ʼ�u�0�&�!�6�}�ϻ�����\l�N��X����2�0�!�8�;�>�������[��v-��Uʜ�u� �;�u�"�}��������P��U�����8�;�1�7�w�����
����c��R!��#���1�0�u�<�?�}�W���T�ƿ�V��V����� ��u�'�$�8����)����|��Y>��ʦ�;�0�&�0�#�<�'�������^F�������3�&�=�&��>�ϼ�Y����P
��\N�����{�u�u�u�$�8����:����P
�
N�����'��9��:�f�W���Yӕ��_��V�� ���9�1�6�u�j�.��������P2��GN��U¦�4�6�=�&��)����-����R�������6�=�&��#�3����7����R��V�� ����%�|�n�]�}�W���TӶ��V
��RN�����4�0� �u�0�4�W���Y����A��������0�3�;�2�����
����U��=N��U���x�<�&�#�;�8��������[��T�����u�;�!�&�4�8��������\	��GN��ʦ�4�!�4�u�2�2�}���Y���2�������0�&�4�0�w�8�϶�����Z��C�����,�&�9�!�>�:��������_��X �����u�u�x�u��1�'�������Z����U���!�{�u�u�w�.��������F��[N�U���4�0�6� �l�}�W���
����c��R!��9���<�0�i�u��1�'�������P
��y������!�x�u�8�3�ϵ�����@��C��6����4�0� ��1�������N��X�����3��1�-�8�	����:����]��Y�����&�&�4�6�?�.�8�������]��������0�3�;�2�����
����_��C��\�ߊu�u�u�x��1�Ϫ�Ӕ��GF����U���%�!�u�;�w�$����Ӌ��P��_�����<�0�1�9�.�4�}���Y�����T����� ��9�<�2�W�W���Y����G��t��9���<�0�i�u��.��������_]ǻN��U���9��4�0�"���������VF������4�0� ��;�9���Y����]��QUךU���u�'�6�&�l�W�W��8����]F��RN�����&�u�&�0�#�<�'�������R
��R�����!�4��4�2�(�!�������9F��y��8���=�&��!�k�}�9���4����R��B���ߊu��&�4�#�<���Y����G��t��9���<�0�_�u��1�'�������R
��R�����6�=�&��#�<��������l�D-�����&��!�i�w���������G*��g��N���;�u��n�