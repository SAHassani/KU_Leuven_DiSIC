-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B"��e�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������4ǶN����d�u�4�u�g�n�Z�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���6�u�e�f��-����Ө��Z	��[N�����8�;�&��%�2�������r
��e�����0�0�#�1�z�}��������]��B�����;�0�;�9��;������ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�x�u�?�.����������C�����&�4���o�}�Ϭ�����]��V�����'�&�9�u�6�6��ԑTӒ����@N�����1�8�<�{��}�Ϻ�
����WF�������4�<�9�u�>�5�!��/��ƴF��SN�����u�{�x�_�z�	�Ϲ�����@F��V�����;�u��!�"�
��������VF��R
��ʦ�0�<�,�"�2�8����T�ƾ�F��PN�����{�u�r�0�8�1�W�������[��@��U���&�u�:�7�9�)����s��ƴF��C��O���z�y�m�d�w�.����U����Q��N�U���0�0�u�<�$�W�Zώ�Y���F�B�Y��}�<�;�1�w�l����U����Z��P�����|�x�u��;����Y����V��^��3���_�x�>� �'�)����Y���]Ƕd�U���u�:�0�u�`�?�����Ʈ�Z��E�����:�3�"�!�w�}����Ӊ��D��DL�����;�{�x�u�?�.��������_��R
��ʦ�!�<�2���6����
�Ƹ���^��E����_�x��s�Y��Y������I�\ʴ�1�&�!�<�0�)�Ͻ�����]F�������}�b�{�x�]�p�>����ƾ�F��X�����<�;�h�e�b�}��������F��EN��U���<�<�0�u�?�}����ӏ��K��X�����%�u�=�;�#�8�W�������@F��P�����=�u�0� �#�4�W�������W	��N�����x�u�<�9�:�4����Y�ƶ�A	��^�����&�2�4�&�#�<�W���Y����R��M��U���&�1�u��>�W�Zϩ�����\��R����:� �0�4�!�/�W����ƫ�Z��E��[���3�,� �'�w�3�Ϭ�����Tl���U���0�u�<�&�w�2�W�������@��_�����1�=�9�u�!�3�W���5����v1��Y�����x�u� �u�1�$�Ȭ�Y����W����U���,�7�!�u�2�:�W���PӒ��]F��RN�����=�:�u�3�z�}��������F��uN�����,�2�0�u�6�}����Y����G��P��U���:�u�%�'�6�5���s������C�����u�:�;�<�0�2���Y����F��SN��ʲ�<�u�'�:�w�<�W������F��_�����"�&�4�:�#�l�;����ƫ�Z��E��U���'�u�e�y�g�}����
���9K�gN�U������u�z�	����
ӑ��GF�������1�<�u�:�2�8�}��T�Ɯ�[��,��U���u����]�p�6՜�E�Ƨ�R
��D�����'�6�<�%�#�W�Zϝ�E�ƈ�G��=C�6�����i�u��)�>���N���9K�c��ʼ�u�u�%�6�6�}����UӅ��z��B��Yʢ�<�=�6�;�2�)�W���������C��4���_�x�<�%�#�2�W���Y����H�c��U��� �u�&�r�w�.�Ϸ�
����G��s=��M���!�&�;�!�>�W�ZϪ�Ӄ��R��YN�����4�:�0�y�?�*��������Z��B
��U���!�0�%�'�w�<�W�������9K�C��U���a�u�:�7�w�1��������G
��Y��U���!�0�%�0�>�(�W���M���`��RN�����u�� �u�i��>�������G����U���,�:�6�'�8�}��������`6������u�&�4�x�w�2��������R��XN�����u�=�u�:�9�8�W���^�Ƽ�R�������:�%�&�!�w�4�ϱ�s����[��g)�����;�u�s�{�w�8�����ƅ�vF��SN�����_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T����Z��E�����_�u�&�u�2�8��������lW��@���ߊu�&�u�0�2�3����������dחXʦ�;�=�&�&�#�<��������9*��E��U���<�-�:�0�>�f��������}/��zU���������8�-����
ݧ��l������<�u�'�;�;�)�(���s����Z��r�����;�0�u�&�w�:�������F��V�����u�!�
�:�>���������W	��C��\��u�w�e�e�g�m�1���B�����C��"���=�o�<�!�0�/�M���H����F��E��U����>�u�u�w�}�MϷ�Y����_	��TUךU����!��u�w�}�W���
����\��h�����a�u�:�;�8�m�L���YӅ��z��B��U���;�&�1�9�0�>����������Y��E��u�u�6�;�"�-����Cӏ��@��[���ߊu�u��!��)�W���Y����@��[�����6�:�}��#�(� �������\��XN�U��0�1���'�2����B����A��C�� �����:�u�&�.�%�������@lǻ�����;�u�&�a�2�}�WϹ�����l�N��4�����u�u�w�}�W���Y����T��S��N���u�u�� ���2���Y���F��^ �����o�u�n�u�w�}�6���Y���F�N��U��<�!�2�'�m�}�L���Y����f2��r=��*�����
���	�W���Y����Q	��R��O�����n�u�w�}�6���+����l6��c+��*��������}�W������F��v:��W�ߊu�u�u�
���W���Y���F������o�u�����}���Y�Ǝ�r5��r)��U���u�u�u�u�9�8����D����F�N��0���u�u�u�u�w�}�W�������AF��_�U���u�����}�W���Y���	F��E��U��w����l�}�W���:����z(��pN��U���u�o�<�!�0�/�M���B���F��v<��<�����u�u�w�g�������F��=N��U�����u�u�w�}�W���Y����]��R��H��_�u�u�u���W���Y���F�T�����0�!�'�o�w��1���?����u �=N��U�����u�u�w�}�W���Y����]��R��H��_�u�u�u��	�6���0����F�T�����0�u�h�d�]�}�W���)����a#��N��U���u�u�;�0�2�}�J��s���F��c:��;���u�u�u�u�w�}��������\�oL�E��e�e�e�w�]�}�W���+���F�N��U���u�u�;�0�2�}�J��s���F��{1��&���u�u�u�u�w�}�������+��|L�U���u������9���Y���	F��E��U��w����u�W�W���Y����a)��s'��*����u�u�!�>�:�M���*����r5��d��U�������w�}�W���Y����@��Y	��H�����n�u�w�}�"���4����F�N��U��&�'�;�u�j��"���*��ƹF�;��*�����
���	�Mϭ�����	[�y!��4����n�u�u�w��2���4���F�N��Oʦ�'�;�u�h�u��C���B�����CFךU���u��u�u�w�}�W���Cӏ����h�����_�u�u�u�w�}�W���Y���\��YN�����:�<�
�0�#�/�E�������V�=N��U�����u�u�w�}�W������G��X	��*���!�'�g�u�8�3���B���F��t!��U���u�u�u�o�8�)��������l��C��G���:�;�:�e�l�}�W���;���F�N��U��<�u�&�1�;�:��������Q��X����n�u�u�u���W���Y���F��^ �����9�2�6�#�4�2�_������\F��d��U������u�w�}�W���Y����@��[�����6�:�}�b�3�*����P���F�tN��U���u�u�u�u�w�3�W���&����P9��T��]��1�"�!�u�~�W�W���Y���F�N��U���u� �u�!��2��������R��S�����|�_�u�u�w��9���Y���F���U���
�:�<�
�2�)���Y����G	�UךU���u�� �u�w�}�W���CӉ����h�����0�!�'�a�w�2����I��ƹF�-��'���u�u�u�u�m�4�Wϭ�����T��=N��U�������w�}�W������G��X	��*���!�'�f�1� �)�W���s���F��e<��4����u�u�u�9�}��������l�N��6������ �w�}�W���Y����F
��^�U���u����w�}�W���Y�ƥ�F��S1�����#�6�:�}�w�2����I��ƹF�/��8���u�u�u�u�m�4�Wϭ�����Z��R����1�"�!�u�~�W�W���Y����j/��r"��U���u�;�u�!��2��������T��X����n�u�u�u���$���0���F��^ �����9�2�6�_�w�}�W���-����|3��N��U���u�!�
�9�0�>�}���Y�ƃ�v4��x9��U���u�u� �u�#��������F�b ��'����u�u�u�w�(�W���&����Z��N��Uʅ�������W����ƿ�W9��X	��N���u�u�����2���-����\��D�� ���<�n�u�u�w��6���Y���F�N��Uʦ�1� �:�<�l�}�W���:����F�N��U��<�u�&�1�"�2���Y���%��{;��1���u�u�o�<�w�.��������9F�N��0��u�u�u�u�w�g����
����_	��TUךU���u��g�u�w�}�W���Cӏ����h�����_�u�u�u��}�W���Y���\��YN�����9�2�6�_�w�}�W���8����}F�N��U���u�!�
�9�0�>�}���Y�Ə�p2��N��U���u�u�;�u�#��������F�t+��U���u�u�u�u�w�3�W���&����Z��N��Uʖ�������W����ƿ�W9��X	��N���u�u���w�}�W���Y����Z�D�� ���<�n�u�u�w��#���Y���F�N��Uʦ�1� �:�<�l�}�W���+����%��e7��U��<�u�&�1�"�2���Y���4��v"��:���u�u�o�<�w�.��������9F�N��&���u�u�u�u�w�g����
����_	��TUךU���u���u�w�}�W���Cӏ����h�����_�u�u�u���%���Y���\��YN�����9�2�6�_�w�}�W���4���F�N��U���u�!�
�9�0�>�}���Y�ƞ�g6�N��U���u�u�;�u�#�������ƹ�������;�n�_�u�>�3�Ͻ�����	F��S1�����#�6�:�}�`�9� ���Y���F��C����e�|�_�u�>�3�Ͻ�����]F��D�����6�o�u�e�l�W����s����p��N'��I���:�u��!��u�@��s������T����0�2�;�'�4�0��ԜY�ƭ�R��R	��K��_�u�u�9�:�9����D����9F�����u�y�x�u�?�.����
����Z��R��ʳ�'��'�0�w�}��������UF��R	�����0�u�:�e�w�4�����ƭ�R
��R
�������u�=�"�5����8Ӌ������U����u�=�u�������Ƹ�VF��C�U���4�!�'�&�#�-��������V��
P�����y�u�u�4�#�/����	����A��R�����!�;�u�k�u��4���s���R9��G��H������w�]�}�W���
����[�BךU���'�2�h�u�{�}�Wϼ�����[�*��0���y�u�u�6�%�$����Y���F�N��'����u��_�w�}��������A��
P��Y���u�6�0�u�i�l�W��Y�ƞ�tl�N�����k�-�f����1���[���F��R	��K��_�u�u� �#�<�������F��=N��U���:�0�0�u�i�m�}���Y����V��
P��W��e�e�e�e�g�q�W���	����X�N�U������u�w�.��������T9��D��K����
���{�}�Wϭ�����XF�L��&���_�u�u�0��<����Y���c'��r<��Y���u� �0�8�;�}�I���6���9F���*���!�'�
�0�2�)�J���7����g"��BךU���&�
�<�1�j�}�8���A����\��Z�����u�9�u�k��6�}���Y�����[����u�:�;�:�f�t�}���Y�����[����u�:�;�:�g�q�W������P"��V'�����u�4�'�<�w�c��������9F�����u��� �"�8�[���Yӄ��]F�F�����u�k�r�r�{�}�WϮ����N��_��U��r�r�y�u�w�>��������[�^�����u� �!�<�9�3�J���I��ƹF��T��U��:�0�y�u�w�?����D�ƣ�V�N�����,�4�6� �w�c����U�����C�����u�k�:�0�{�}�WϮ�D�Ư�U��d��Uʥ�!�0�;�1�#�>�W�������9F������1�!�6�u�i�2���Y����E��[��H���%�;�_�u�w�3�������	��YBךU���4�'�:�!�j�}����s���C��CN��U���;�_�u�u�'�2���Y����V��BךU���9�8�1�u�i��G��U�����E�����h�u�e�e�{�}�WϽ����A��d��Uʶ�4�u�k�r�p�W�W�������\��
P��D���u�u�6�7�w�c�P���s���P��S�R��_�u�u�0�w�c��������u �N�����'�,�;�h�w�l�[���YӅ��[�_�����u�0�!�9�j�}�F��Y����V�	N��R�ߊu�u�0� �#�<����Y���A�N�����u�k�r�r�]�}�W�������W�	N��R�ߊu�u�&�7�j�}�G��Y����@��
P��E���u�u�'�!�;�>�������V�=N��U���8�h�u�e�{�}�WϬ�����[�^�����u�&�%�h�w�m�^�ԶY���g��{=��U���0�7�0�u�8�3��������V��C��8���_�u��!��)�K���)����R��S�����m�>� �%�#�4����s����4��d