-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����0�:�,�#�3�p�W�������y	��/�����;�x�u�'�0�3�ώ�����	F��~��C���_�x��!�m�o�W��� ����l�=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z�u�^��H�Ə�C��P��;���:�4�u�;�#�(����Y����\��^��X���9�u�<�=�$��������(��^��ʜ�&�'�8�;�$������ƅ�U	��V�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԑTӶ��C	��N�����3�9�u�'�6�8�W���Y������X�����!�0�3�4�#�2��������G	��=C�U���u�u�u��>�}��������Z��V �����u�u�<�%�2���������a'��V �� ���u�0�1�"�>�8�Z���Y���F�G�����u�:�8�>�w�5�ϳ�����Q��A�����4�#�'�4�;�}����ӕ��U��R	�����_�x�u�u�w�}�Wϊ�Ӌ��\��T�����0�`�g��w�<����W���K�N��U���u�=�u�4�6�4�W���Y����Z��YN�����:�u�<�;�3�e����&�Ʃ�V��C�X���u�u�u�u�w�5�W���������C��4���<�0�4�1�<�<����8����I��R��ʡ�0�x�u�u�w�}�W�������UF��RN�����;��!�%�%�.��������V
�������!�'��/�]�p�W���Y�����R�����!�0�&�0�w�)� ���Ӓ����SN��ʡ�4�0�&�&�#�8������ƴF�N��U���>�4�4� ��$����
����WF��CN��U���2�'�!�4�w�����8����I�CחX���u�u�u�u�$�8��������F��DN��ʧ�4�u�1�'�$�}����
����WF����ʡ�u�=�_�x�w�}�W���Yӈ��GF��X�����u�;�!�_�z�p�W���Y���F��RN�����1�'�&�u�8�3����
Ӊ��JF��S��ʢ�0�u� �1�#���������9K�N��U���u�<�u�'�2�}�#���	����V��DN�����u�<�=�&�2�9����
����D��=C�U���u�u�u�&�8�9��������@/��V�����u�!�0�"�$�}�Ϸ�Y����V��C�����x�u�u�u�w�}�W�������Z��E�����:�!�0�;�/�}���� Ӈ��A����ʦ�4�4�;�4�>�W�Z���Y���F��D����� �0�>�;�%�0����8����Z��EN��U���0�!�<�u�?�}����Y����V��C��U���u�u�u�:�9�8�W�������G��EN�����0�!�u�=�9�.��������W6��RN��U���0�_�x�u�w�}�W���.����X/��E������1�:�;�2�}�Ϫ��Ƹ�VF��Z��U���4�0�u�<�2�<�;���s���F�N��U���:�,�"�!�w�}����������E�����4�1�0�&�w�5�ϵ�����V��E/��%���!�'�x�u�w�}�W���Y����R
����U���:�,�4�!�w�4�Ͽ�?����^��E�X�߇x�u�u�u�w�}��������Z��_�����!�4�u�4�w�8�ϸ��ơ�^	��d����u�u�u�u�w�	�Ϯ�	����VF��[�����u��4��6�����
����]��b�����4��1�0�$�p�W���Y���F��SN�����1�'�&��w�2��������Z������,�9�&�_�z�p�W���Y���F��RN�����;�u�0�4�w�/�ϭ�����R��S�����4�1�&�%�6�8��������@l�N��U���u�u�;�u��<�6���������D<�����'�&��!�>�}�W����Ư�P
��=C�X�߇x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s����R��^��Yʢ�'�n�u� �2�4��������T��_�[���n�u� �0�>�8�Y�������@��V�����&�u�:�>��:��������@"����N��� �0�"�'�y�6�3�������F��RN�����>��4�!�2���������@H��[Uװ���!�u�'�6��>����������N�����6�_�u�u��>��������W6��Y��U��<�u�:�9�6�}�JϪ���ƹF��s��<���,�<�0�u�w�}�W���Y����]��R�����u�u�:�g�w�`�E�ԜY�Ƨ�R��B�����0�u�u�u�w�g��������AF��Y	��Dʡ�u�u�o�u�~�W�W������F��Z��6���o�<�u�!��2���s���@4��R�����1�'�&�u�m�4�W�������9l�N�����0�1�1�'�$��W���ӄ��_��d��Uʦ�%�4�0�0�3�9����Y�ƥ���[��N�ߊu�u�x��2�3����Y����Z��C�����&�u�d�u������
ӂ��V��������!��,�>�8�}���Y����W'��E��<���u�;� �&�0�8�_���K����N��A����� ��,�<�2�}�������K�bV�U��� �{�_�u�w�.��������WF��^ �����4��6�:������8����I�_�����:�e�n�u�w�.��������Z��^	�����'�4�
�}��)�>��� ����K�
�����e�n�x�u�f�s�}���Y����R/��T��ʆ�2�0�d��%�$�ǵ�����r��^��X��1�"�!�u�~�}�Zύ�A��ƓF�D*������o�:�!��:���8����l��s��:���'��/�u�w�}�������K�d_�D���u�&�4�4�"��Mϱ�ӵ��]��/�����}��!��#�/�$���Y����W	��C��\���x��m�d�]�}�W�������A��x��Oʺ�!� �&�2�2�u��������W��\*������,�<�0�w�2����I����K��@����l�l�0�1��<����=����V��NUװ���<�0�!�'�w�	�W���?����w��V�����,�<�_�u�z�}��������Z��T�����&�1�3�;�w�5�W���Ӏ����
�����;�u� �;�>�4�Ϫ����K��R�����u�=�u�<�2�2�W���Y����A��Y�����_�u�:�&�6�)����=����Z��T�����0�u�h�f�w�}�3���0����`��d�����4�u��8�2�9��������]��R����<�;�9�&�6�<��������V'������u�h�3�9�2�W�W�������w��~ �����<�0�u�u�8�1��������X"��V'�����/�x�u�:�9�2�G���D�Σ�[��S����0�n�u�&�0�<�W�������Z��T�����1�m�'�4��u�3���0����`��C��U���;�:�e�u�j�u����
���	��R��H���e�|�n�x�w�l�Y�ԜY����R
��s��<���%��o��0�8�Fן�������C��4���<�0�x�d�3�*����P���	��R��H���:�=�'�u�i�z�P���Y����^�=N�����9�&�0�0� �4��������Z��N�����;�o�u�4�$�f�}���TӲ��$��zN�����!�'�u�d�w�����
������DN��ʥ�<�|�u��>�8����
���F��R
�����2�u�<�&�#�}����
�ƭ���V��ʦ�/�u�d�u�w�����8����Iǻ�����!�>�'�!��9��������\��Y�����h�:�g�`�e�6��������Z��d�����4�u��<�2�9����Y�ƹ�@��R
��"���0�1�'�&��3����Y�ƨ�D��^��O���:�=�'�u�i�z�P��Y����
H��X��M��_�u�x��2�}�3���8����I��DN�U���d�-�g���}�ϫ��Ƹ���G��U���!�;�u�u��.����
���F��R�����0�u�9�=�"�5��������JF��YN�����`�g�g�d�e�}�&ϭ�����F��[��D����u�x�u�6�-�����ƾ�B��R
����!��1�0�$�>�ϼ�Y�ƣ�_��^�����y�u�7�!�#�8�������K��S
�����&�4�"�,�w�}��������'��^ �����<�!�u�<�9�1����
����\F��V�����u�x�u�1�%�.�W�������9F��^	��ʦ�0��<�0�3�/����Y����T��V�����:�e�u�h��)����D���O��C� ���_�u�&�2�6�}�%���8����@������1�&�0�1�3�/����^����VO��F�����u�k�r�r�l�}�����ƿ�V��S
�����;�&�;�u�w�3����ە��R��S�����'�;�0�n�]�}�Z���Ӓ����VN��U���4�u�&�2�2�)�Ϫ��Ƹ�VF��C�� ���!�0�8�8�%�}��������@l�C�����u�;�u�=�;�2����Ӈ��\��S��U���u�4�4�9�;�.����ӑ��G��'�����u�4�0�u�z�}��������@��^�����7�!�u�3�#�8����Y����V��G�����7�6�8�u�9�2����WӲ��9F�N�����u�4�u�0�"�8�W���
����GF��^�����<�;�3�:�w�5�W���Ӆ��Z��X�����=�_�u�x�:�0��������G	��s��:���_�u�:�&�6�)����6����G*��P��Oʼ�!�2�'�o�w�2�Eǵ�����r��^��Zʾ�4�4� ��.�4���Y���g��[�����d�|�3�;�#�2�W����ƾ�G��DN�����#�u� �7�%�s����
ӕ��V��_��U���u��8�3�$�)��������\F��Q��U���2�&�_�u�8�.��������U ��C&����<�!�2�'�m�}��������X"��V'�����/�u�u��#�����*����l�D������8�3�&�#�g��������X+��x�����2�u�:�;�8�m�W��Q����A�	N��R��u�&�2�4�w�����
����C��N�����0�}��8�1�.����ӂ��]��G�Uº�=�'�u�k�p�z�L���
����_F��R������%�d�o�"�.����Q����| ��R�����:�;�:�e�m�}�������A��UךU���;�9�&�0��<�6��������^	����1�"�!�u�~�g�WǱ�����X�I����,�0��#�a�/����Y����A�� �� ���u�4�2�i�~�2�W���&����P9��T��]���1�"�!�u�~�W�W�������~��V�� ���o��2�0�f�����ۍ��G��v�����x�d�1�"�#�}�^���Tӵ��W��\ךU���;�9�&�0��)�8���Y�Ɵ�T��V�����!�>�4�4�9�/�$���Y����W	��C��\���x��m�d�/�o�}���Tө��C��^ �����/�!�:�_�w�4����
����|��{��Oʆ�2�0�d��%�$�ǵ�����G'��d��U���u�:�;�:�g�}�J�������[������h�u�e�|�l�p�W��W���@��V��1����!��9�m�����H˧��R�������!�'��/�w�}�W������F��F�����u�k�}�!�2�.�J���I���K�d_�D�ߊu�!�'�7�#�}����Cӕ��Z��=N��Xʐ�&�'�u�=�#�)����
����_��E�����0�2�1�"�#�}����Y����@	��_�����'� �<�2�3�1����T�Ƹ��������<�u�=�'�]�}��������X�������0��<�0�3�/����	����Z��[N��Uȡ� �w�_�u�#�/����Y����	��D#��'����1�0�&�w�4��������A��d�����<� �0�>�2�}�ϭ�����e��S>����&�2�4�u�$�����B����G��U��U���%�:�u��#��!�������q\��^	��ʼ�u�!� �w�]�}��������X�������4�;�<�0�m�.����Y���G��UךU���'�7�!�u�2�-����=����]6��R?����4�u�&�w�%�8�L�������Q����ʺ�u��!��#���������������u�4�!�<�"�8����Y����w��x��9���u�<�;�9�>�}����[��ƹK��_��*���&�4�!�u�z�+����
����Wl��R	�����x��%�9�9�}����=����]0��^
�����9�&�u�=�$��W���Y����_��SN�����!�u�=�u�2�2��ԜY����G��@��U���u�:�!�;�w�8����Ӓ����X�����1�6� �0�6�)����Y����F��=N��Xʛ�!�u�=�!� �}��������]��@�����&�:�u�=�$�)�W�������R��BךU���6�&�}�4�'�8����Yӄ��ZǻN��ʧ�&�;�
�1�2�����:���G��=N��U���x��<�u�>�8����Y����WF��R��ʼ�6�0�0�!�#�8� ���Ӈ��A�������_�u�u�u�z�*�����Ơ�@��[�����;�!�0��#�}�Ͽ�����@F��[�����u�u��!����������[��s��<���9�1�>�4�6�3�������O��=N��U���x�=�&�%�'�1����������DN��U���u��!�'�>�<�W�������V��N@ךU���u��!���1���������C��#���1�_�u�u�9�}��ԜY����C��R�����x�u�<�0�>�8����
����z��^	��ʦ�u�=�&�u��}����Ӗ��P��T��ʡ�u�=�u�0�8�$�}���TӉ��V��D�����:�!�;�u�2�<�W�������V��NN�� ���6� �0�4�#�0��������VHǻ�����}�4�%�0�;�t�Wϼ���ƹF��QN�����
�1�0��:�1�4���Y����9F�N��1�����%��k�}�3���0����F�N�����;�<�0�u�j�.������ƹF��Y
���ߊu�;�u�'�4�.�L�ԜY�ˏ�V����U���!�u�1�'�$�}�������C��R��&���9��>�_�w�8��ԜY�ƥ���^ �����}�4�%�0�;�t����s���F��R��"���0�1�'�&��-�W��
����G1��C�����&�_�u�u�w�;��������G��S�����0�!�0�_�w�}�W���.����r��R��I���:�=�'�u�i�z�P��Y�����^��1�����9�1�>�8�^Ϫ����F�N��U���6�0�0�!�%�9�'�������[��N��U���u�&�'�!��9����E�ƿ�A��v
�����~�d�_�u�w�}�W������F�N��"���0�1�'�&�w�`��������A��C��N���u�u�u�0�3�4�L���Y����]��QUךU���;�u�3�_�w�3�W�������9l�C�����;�&�'�!��9����ӕ��^1��C�����&�u�3�&�2�
��������@F�������0�4�9�_�w�p����I�Ƹ�VF��U@ךU���6�&�}��>�8����
��ƹ��^ ךU����8�'�!��9����E����G��DN��U��|�_�u�u��0����8����@��`�����'�&�r�4�0�t�K���.����r��R�����;�u�'�6�$�f�}���Tӥ��R��C��'���u�1�'�&�w�2����s�Ƽ�\��DF������>�_�u�2�4�}���Y����Z��P1�����4�%�0�9�~�)��ԜY���Z ��b�����4��1�0�$�)��ԜY���F�������4��1�0�$�3�W������F�N��'����1�0�&�k�}�%���8����@��d��U���u�0�&�_�w�}�W���Y����W'��E��U��&�0�1�1�%�.�:���
����9F�N��U���u�3�_�u�w�}�������F��SN��N���0�1�%�:�2�.�}���
����r��R������0�i�u��<�6������W��=N��Xʅ�%�9�;�u�?�}�%���8����@��^	��ʦ�u�=�&�u��}����Ӗ��P��T��ʡ�u�=�u�0�8�$�}���TӉ��V��D�����:�!�;�u�2�<�W�������V��NN�� ���6� �0�4�#�0��������VHǻ�����}�4�%�0�;�t�Wϼ���ƹF��QN�����
�1�0��:�1�4���Y����9F�N��Xʜ�u�=�u�4�6�3���� ӏ��_��R�����!�0��!��)�W���Y����A��Y�����!�1�=�&�w�}�W��Y�ƨ�G��B�����<�u�0�0�6�}�&ϭ�������R@������u�3�&�2�9����
�ƭ�Vl�N��X���&�1�1�'�4�1�W�������~��R�����&�{��0��?� ���Y����@��C�����!�!�0�u�w�}�Z�������WF�������:�u�u�4�6�2�ϓ�!���F�D#��'����1�0�&�k�}�������A��U��Xʱ�3� �!�4�$�:����W���F��z�����1�'�&�}��<�6�������Z��N�����3�0��;�#�}�������[��e��4���0�&�&�0�3�9����^������Y������3�0��9�)�^�ԜY�Ʃ�WF��d�����%�:�0�&�]�}�Z�������GF��RN�����_�u�x��:�1�W���Ӷ��GF��zN��1���<�u�=�u�8�)����������[�����<�;�3�'�#�8����Y����A��dךU���=�:�
�u�%�>�3�������CF��V�����x�#�:�>�0�6��������VF��V������/�_�u�z�5����Y����G��S��ʦ�0��<�0�3�/��ԜY�˺�\	��VN�����;�4�<�u��)�>�������C��N����>�4�&�4�6�3�W�������Z��=N��X���:�
�u��#��&ϭ�����c��fd��Xǣ�:�>�4�&�2�9����
�ƿ�V��V
�����&�u�x�#�8�6�ϭ�����G/��z����� ��u�x�!�2����
����|�������4� ��u��<�$���Y����G��X��3���!�0��4��-�_���P�����R��U���u�_�u�u�w����� ����[�\*�����'��/�|�w�p��������V��V ��U���:�g�o�u�]�}�W���Ӌ��NǻN��U���%�0�9�u�w�}�Iύ�����_�N��U���u�x�<�u�$�9�������F��`�����'�&�u�k�$�8� �������V��N��Xʼ�u� �&�2�2�u�W������l�N�����4�;�4�<�w�`�W�������R
��g��7���x�u�;�u�8�1��������X"��V/��&���x�u�:�;�8�m�}���Y�ƿ�R��Y'��U���h�u��!������Y���F���U���;�1�m�'�6��_�������`��_�����:�e�u�u�w�.�������F�	N�����;�<�0�y�w�}�W��Y���`��R
�4���,�!�>�4�6�/�$���T�ƨ�D��^ךU���u��4��3�8����Gӕ��^4��S/�����y�u�u�x�>�}��������F��@ ��U���u�u�u�&�6�<����Y���F��R�����!�y�u�u�w�p�W���Y����V��v�����>�4�4�'��'�Z�������VǻN��U���!��!�u�w�}�Iϭ�����R)��fG�U���u�x�:�!��:���8����l��s��4���<�0�d�1� �)�W�ԶY���@+��s��:���z�u�&�1�;�$�������@F��C�����6�u�:�!�2�.��������@l�G������8�9��<�W�W������F�������0�2�}�4�'�8��������F�N�����3�0�u�h�$�8��������X+��x�����2�u�:�;�8�m�L���Y����~��Q�����0�u�h�&�2�����B���F��z�����!�<�0�u�j�.��������Z��d��Uʰ�1�<�n�u�2�9��������9F�N�����u�u�<�;�;�)�W���������C��U���!�0��8�%�}����=����1��YN�����;�'��/�]�}�ZϷ�Y����G��C��U���!��!�'��'�W�������V��G����!�u�:�!�2��W���	����\ ǻC����'�&�u�<�?�3����=����r��N@��ʡ�0�u�'�u�&�<�W���ӈ��\ ��R��ʻ�0�0�u�;�]�}�Zϭ�����@��^��U���;�!� �0�y�}����+����U ��CN�U���=�;�>�0��;��������F��R��U���<�!�2�'�$�8�8�������VW�=d��X��� �u�;�u�>�8��������R��X�� ���:�8�>�u�>�4�ϻ�
�Ƹ���CN�����;�!�0�8�:�/�}���TӇ����#��[�ߊu�x��9�4�}����������C�����!�:�3�0�y�}�0�������G'��d�����<�<�u��#�����*����F��S�����u�0�0�4�2�}�WϮ�����5��G�����u�u�7�2�9�}�W����ƾ�@��h���8�9��>�w�5����Y���F��s��:����9�<�u�j�.��������zN��R�����3�0�u�u�~�W�W���Y���@"��V!��$���}�|�i�u��0��������~��R�����!�~�<�n�w�}�Wϻ�ӏ��9F���U���6�&�n�u�2�9��������t��V�� ���,�_�u�x�w�.��������F��CךU���!��!�u�j�.��������_]ǻ�����!�u�h�&�6�<������ƹ��V
�����&� �u�h�$�8��������Z��x �����u��n�