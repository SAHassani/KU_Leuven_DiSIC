-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B"��V���߇x��!�:�m��Ϝ���ƴF��^	�����'�?�6�o���(��L���"��RT��Bʟ�;�4�,�g�f�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�CחX���|�g�d�u�8�$����Y����\��'�����0�!�u�:�'�/����s����_
��^	��ʇ�&�'�0�_�z������ƅ�@��Z��ʜ�!�'�4�u�9�2�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�x��>�}��������Z��V �����u�u��a�{�>��������U	��VN��6ʺ�u�6� � �6�8�}������Z	��N��U���1�&�;�0�w�2��������Z����ʃ�y��y�4�3�����Y��ƴF�N��R���;��x�u�w�}�1ϱ�Y���F�(�����u�x�u�u�w�8�}��YӶ��VǶN��Dʓ�u�;�:�8�3�W�Z��Y�Ƨ�P��B�����4�&�_�x�w�}�'������F��uE�����:�8�1�h�g�l�F��s�����T�����'�!� �_�z�}�Wώ�)����Z�N�����u�=�;�6�4�(��������F��Z��H��d�d�e�_�z�}�Wώ�)����Z�gE�����u�=�;�6�4�(��������F��Z��H��d�d�e�_�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǑ=�����u�0�0�_�w�.�W���ݕ��l
��^��D��4�9�_�u�$�}��������Z��C
����_�x�&�;�?�.�Ϫ�����G��Q�����'�u�<�<�/�2����B����A��;��&���_�&�u����!���	����G��{"�X���,�!�0�<�w�/��������9l��Y��ʐ��%�m�<�w�W�W�������9F������;�=�<�u�w�}�ϼ�����\�Q���ߊu�u��6�:�1����Y����Z��X�����h�3�9�0�~�W�W������F��\N��Oʼ�u�!�
�:�>�f�W������\��YN�����2�6�#�6�8�u�@Ϻ�����O��N�����d�o�<�u�#�����B�����v\��U���&�1�9�2�4�W�W���;���	F����*���<�
�0�!�%�l�W������]ǻN��0���u�u�;�&�3�1����s���P6�N����&�1�9�2�4�+����Q����\��XN�N���u�6�;�u�m�4�W���&����P]ǻN��%���u�u�;�&�3�1��������AN��
�����e�n�u�u�4�>����Y����@��[�����6�:�}�b�3�*����P���F��T!��U��� �u�!�
�8�4�(������
F��@ ��U���_�u�u��4�0����Y�ƥ���h�����n�0�1���-�O�Զs����Z��C��U���u�3���'�e��ԶYӅ��C	��Y����0�u�u�2�9�/��ԜY���r%��t<��U���u�u�u�u�w�3����Y���l�N��4������u�w�}�W���Y����T��S��N���u�u���w�}�W���Y���F��^ �����o�u�n�u�w�}�6���+����l6��c+��*�����u�u�w�}�W�������	[��v"��N���u�u�����#���-����l"��r-��:����u�u�!�>�:�M���4����]ǻN��U���� �u�u�w�}�W���Cӕ��Z��S��1����w�_�u�w�}�4���+���F�N��U���;�0�0�u�j�l�}���Y�Ǝ�v!�N��U���u�u�u�u�9�8����D����F�N��<����u�u�u�w�}�W�������\�*��0���n�u�u�u���.���<���F�N����2�'�o�u�l�}�W���:����z(��{<��U���u�o�<�!�0�/�M���B���F��e+��U���u�u�u�u�w�g�������F��=N��U�����u�u�w�}�W���Y����Z��R����u�w�����1���B���F��e+��U���u�u�u�u�w�g�������F��=N��U��� ������0���Y����]��R��H��_�u�u�u���2���Y���F�T�����0�u�h�d�]�}�W���8����}F�N��U���u�u�<�
�2�)���Y����V��^�E���_�u�u�u���W���Y���F�T�����0�u�h�d�]�}�W���<����`-�N��U���u�u�!�<�0�g�W͓�*����F�N��9������u�w�}�W�������\�>��!���w�_�u�u�w��(���7����l+��|N��U���<�2�o�u���:���[���F�d'��8���u�u�u�u�w�}�W������F��v(��N���u�u� ����W���Y���F��D�����h�w� ���f�W���Yӳ��l6��c+��*�����o�&�%�3�W��[����r2��cL�U���u� ����}�W���Y���	F��E��U��w��a�w�l�}�WϮ���ƹF�-��U���u�u�u�u�m�4�Wϭ�����T��=N��U���u�u�u�u�w�}�W������G��X	��*���!�'�g�u�8�3���B���F��t'��U���u�u�u�o�>�}��������l��C��G���:�;�:�e�l�}�W���8����F�N��U��:�!�&�1�;�:��������_��X����n�u�u�u��}�W���Y���F��^ �����9�2�6�#�4�2�_������\F��d��U�����u�u�w�}�W���Y���@��[�����6�:�}�b�3�*����P���F�u-��!���u�u�u�u�w�(�W���&����P9��T��]��1�"�!�u�~�W�W���Y���F�N��U���u�;�u�!��2��������R��S�����|�_�u�u�w�}�W���Y���F���U���
�:�<�
�2�)���Y����G	�UךU���u���u�w�}�W���Cӏ����h�����0�!�'�a�w�2����I��ƹF�>�� ���u�u�u�u�m�2�ϭ�����Z��R����u�:�;�:�g�f�W���Yӥ��a?��N��U���o�<�u�&�3�(����B���F��v<��:���u�u�u�o�8�)��������l��C��Fʱ�"�!�u�|�]�}�W���8����r5��yN��U���;�u�!�
�;�:��ԜY���p'��n-��6���u�u�u� �w�)�(�������F�N��8���u�u�u�u�w�}��������T��A�����u�:�;�:�g�f�W���Yӧ��~)��N��U���o�<�u�&�3�1��������AN��S�����|�_�u�u�w��%���*���F���U���
�:�<�
�2�)�������\F��d��U��������}�W���Y����G��[���ߊu�u�u� ���9���Y���	����*���2�6�_�u�w�}�!���5���F�T�� ���!�
�9�2�4�W�W���Y����a ��`N��U���u� �u�!��1����s���F��c:��;�����u�u�"�}��������l�N��%��������}�W���Y����F
��^�U���u���u�w�}�W���Y�ƥ�F��S1�����n�u�u�u���W���Y���F��^ ����� �:�<�n�w�}�Wϝ�8����w#�N��Oʼ�u�&�1� �8�4�L���Y����v$��N��U���u�o�<�u�$�9������ƹF�-��G���u�u�u�u�m�4�Wϭ�����T��=N��U����u�u�u�w�}�W������G��[���ߊu�u�u����>���Y�������*���2�6�_�u�w�}�2���5���F�T�����!�
�9�2�4�W�W���Y����F�N��U���u�;�u�!��1����s���F��z;��6�����u�u�9�}��������l�N��6���u�u�u�u�w�}�W���Y����F
��^�U���u���u�w�}�W���Y�ƥ�F��S1�����n�u�u�u��	�;���+����F��^ ����� �:�<�n�w�}�Wό�-����|"��N��Oʼ�u�&�1� �8�4�L���Y����`2��N��U���u�o�<�u�$�9������ƹF�<��6���u�u�u�u�m�4�Wϭ�����T��=N��U������u�w�}�W������G��[���ߊu�u�u���}�W���Y�������*���2�6�_�u�w�}�$���Y���F�T�����!�
�9�2�4�f�Wϻ�Ӆ��C	��Y����<�;�9�6�2�)�W��
����\��h�����g�u�:�;�8�m�W��Q����A�^��N���&�2�4�u������Y����_	��T1�����}�u�:�;�8�m�W��Yۉ��V��	I�\�ߠ7�2�;�_�w�����Dӕ��l
��^�����'�'�&�/��4�������O�=N��:���1�u�h�w�g�m�G�������X ��D��6���;�0�&�u�w�p�W�������P��@��U���&�u�;�6�6�3�W���Y���F�^�E��w�"�0�u�8�}�6�������\��[��X���:�8�9���}�W���Y���F�_�D���"�0�u��4�0����D���V
��L�D��e�n�x�u�4�(������ƹ��V����1�%�m�_�w�8����Y����9F������2�h�u�y�w�}��������TF�_�U���4�0�u�k�e�W�W�������@��G�����1�!�6�u�i�;����s���R��E�����!�0�;�1�#�>�(������F��v:��W�ߊu�u�
�;�"�}�I���0����JǻN�����'�2�h�u�{�}�Wϼ����W�N�����%�!�h�u���4���s���P��N�����k�d�_�u�w�<����
����TF�_�U���6�0�u�k�g�W�W������F��(��3�����w�_�w�}����D����9F������'�<�'�2�j�}�[���YӉ��\��R	��K��_�u�u�4�#�/�W�������V��^�E���u�u�%�0�w�c�F�ԜY�ƿ�_9��B �����4�>�h�u���:���[���F��[1�����k�w���{�}�Wϭ�����G��S�W�����w�_�w�}�������F��b"��&���u�u� �0�'�)��������GF�L��*�����y�u�w�(�������D��rZ�\��'�u�4�}�w�}����D�Ư�XJǻN��U��6�0�!�_�w�}�W�����ƹF��S�]���0�&�h�u�g�t�}���Y����J��
P��E���u�u�4�<�w�c�_������F�G�U���7�<�u�k��)����D���O�N�����u�k�6�6�9�W�W�������R��YN��U��y�u�u�8�;�.����Y���A�N�����!�h�u���)�}���Y����GF����ߊu�u�4�'�4�.����D�ƣ�V�N�����&�2�:�!�j�}����s���CF������u�4�!�'�5�8����D�ƣ�V�N�����0�;�0�0�#�`�W������F��R�����k�:�0�y�w�}��������[�X��Y���u�6�'�,�"�}�Iϱ���ƹF��T��U��6�6� �y�w�}���������z��Y���u�4� �:�2�`�W��I����F�T�����0�u�k�w�g��}���Y����[�T+��D�ߊu�u�0�g�j�}�2���U�����[�����k�r�r�_�w�}���D���JǻN����h�u�d�y�w�}����D���JǻN�����'�<�u�k�p�z�}���Y����X��r �����u�0�!�9�j�}�F��Y����V�	N�����u�u�6�8�;�>�������W�=N��U���4�h�u�e�{�}�WϬ�����\��
P��E���u�u�'�!�w�c�P���s���A��S�R��_�u�u�&�6�1�������A��d��Uʧ�!�u�k�r�p�W�W���
����_F�I�Y���u�'�!�u�i�z�P��Y��ƓV��e:��