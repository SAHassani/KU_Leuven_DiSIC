-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��V�����%�:�3�<�>�3�������r��X�?���u�8�0�8�9�<�ϔ�
�Ə�]��Xd�U���2�;�9��8�8����!����R��=C�1���o�e�u� �2�o�F�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�}�|�g�f�}��������}��X ��U���!� �0�!�w�2��������K��[�����&��&�'�2�W�Zϐ�����_F��D�����&��!�'�6�}��������]l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z���������[��Q��U���!�<�&�!�2�>��������@F��EN�����%�&�u�<�#�/��������9K�N��U���u�<�u�u�8�-��������*��a'��[�߇x�u�u�u�w�}�#�������U	��C�����,�6�;�4�9�3�W���Y����U��R ��U����#�c�'��W�Z���Y���F��Y
��ʱ�3�;�1�<�w�5�ϸ�����[�N�����3�0�6�u�;�0����Ӓ����VחX���u�u�u�u�?�.����	����	��^ �����<�;�u�=�w�l����Y����Z ��V �����u�0�'�&�9�W�Z���Y���F��_�����<�<�;�u�#�8����K��������U���9�&�u�<�9�;����Y������=C�U���u�u�u�4�3�1����H���F����U���9�"�;�u�8�;������ƴF�N��U���x�u�u�u�w�}�W�������u��C'�����:�3�<�<�9�.��������G��C�����3�6�0�!�w�3����s���F�N��U���0�4�1�'�'�<��������V��R �����8�u�4�&�]�p�W���Y���6��Q��ʙ�6�!�:�u�1�
��������P��C��6���3�6�0�!�y�4�}��Y���F�N��[���:�'�0��:�2����V����G��V�����:�4�:�z���}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d�����'�u���]�}����<����G��X	��*��a�4�9�_��>����)����R��Y�����3�<�<�;�$�4�}�������`
��/��*���&�4�'�,�w�<����Y����VF�G��ʦ�1�9�2�6�!�>����Lӂ��]��G����:�&�4�!�<�<��������R�=��Fܔ�,�!�f�l�w�2����I���F�N��X����&��0�1�/���Y���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��d�d�d�d�f�l�G��I���F�^�E��e�e�e�e�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��d�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�F��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�d�g�l�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�E��e�d�d�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��e�e�d�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����W��^�E��e�e�d�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��H���F�^�E��e�e�e�e�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�d�d�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�l�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�f�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��d�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�l�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�d�u�}�W���[����W��_�D��d�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��H����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��d�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�F���Y���D��_�D��d�d�d�e�g�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�F��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�d�u�}�W���[����W��_�D��d�d�e�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�F��H����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�e�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��d�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�F���Y���D��_�D��d�d�d�e�f�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�e�e�y�]�}�W��H����W��_�E��d�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�d�u�}�W���[����W��_�D��e�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��I����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�l�[�ԜY���W��_�D��d�d�d�d�g�m�G��I����W�d��U���d�d�d�d�f�l�F��H����V��^�E��d�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�F���Y���D��_�D��d�d�e�d�g�l�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�e�y�]�}�W��H����W��_�D��d�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�l�G��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�d�u�}�W���[����W��_�D��e�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��H����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�d�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��d�w�u�u�w��F��H����W��^�D��e�e�e�e�g�m�F���Y���D��_�D��d�d�e�d�g�m�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�e�e�y�]�}�W��H����W��_�E��d�e�e�e�g�m�G��I���F�_�D��d�d�d�d�g�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�d�u�}�W���[����W��_�D��d�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�l�[�ԜY���W��_�D��d�e�d�e�g�m�G��I����W�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�e�g�m�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�d�y�]�}�W��H����W��_�E��e�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�D��e�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��H����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�e�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�e�g�m�F��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�d�y�]�}�W��H����W��_�E��d�d�d�d�f�l�F��H���F�_�D��d�d�d�d�g�l�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�D��e�d�e�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�F��I����W��_�D��y�_�u�u�f�l�F��H����V��^�D��d�d�d�d�f�m�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��I����W��_�D��d�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�e�d�g�l�F��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�d�d�y�]�}�W��H����W��_�D��e�d�d�d�f�l�F��H���F�_�D��d�d�d�d�f�m�G��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��d�d�d�e�u�}�W���[����W��_�D��e�e�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��H����W��_�D��y�_�u�u�f�l�F��H����V��^�D��d�d�d�d�f�m�[�ԜY���W��_�D��d�d�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��H����W��_�D��e�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�d�e�f�l�F��H����W��L����u�d�d�d�f�l�F��H����V��_�D��d�e�d�y�]�}�W��H����W��_�E��d�d�d�d�f�l�F��H���F�_�D��d�d�d�d�g�m�G��H����W��^�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�D��e�e�e�d�f�l�F��H����FǻN��D��d�d�d�d�f�l�G��I����W��_�E��y�_�u�u�f�l�F��H����W��_�D��d�d�d�d�g�m�[�ԜY���W��_�D��d�d�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��H����W��_�D��e�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�G���Y���D��^�E��e�e�e�e�f�l�F��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�e�d�y�]�}�W��I����V��^�E��e�d�d�d�f�l�F��H���F�^�E��e�e�e�e�g�l�G��H����W��^�W���u�u�w�e�g�m�G��I����V��_�D��d�d�d�e�u�}�W���[����V��^�E��e�d�e�d�f�l�F��H����FǻN��E��e�e�e�e�g�m�F��I����W��_�E��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�g�m�[�ԜY���V��^�E��e�e�e�e�f�l�F��H����V�d��U���e�e�e�e�g�m�G��H����W��_�D��e�w�u�u�w��G��I����V��^�D��d�d�d�d�f�l�G���Y���D��^�E��e�e�d�d�f�m�F��H����W��L����u�e�e�e�g�m�G��H����W��_�D��d�e�e�y�]�}�W��I����V��^�D��e�d�d�d�f�l�F��H���F�^�E��e�e�e�e�f�m�F��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�d�e�d�u�}�W���[����V��^�E��e�e�e�d�f�l�F��I����FǻN��E��e�e�e�e�g�m�F��I����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�d�e�d�f�l�F��H����W�d��U���e�e�e�e�g�m�F��H����W��_�D��d�w�u�u�w��G��I����V��_�D��d�d�d�d�f�m�F���Y���D��^�E��e�e�e�d�f�l�F��H����V��L����u�e�e�e�g�m�G��H����V��_�D��d�d�d�y�]�}�W��I����V��^�E��d�d�d�d�f�l�F��H���F�^�E��e�e�e�d�g�l�G��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�d�e�d�u�}�W���[����V��^�E��e�e�d�d�f�l�F��I����FǻN��E��e�e�e�e�g�l�F��I����W��_�D��y�_�u�u�g�m�G��I����W��^�D��d�d�d�d�f�l�[�ԜY���V��^�E��e�e�e�d�f�l�F��H����W�d��U���e�e�e�e�g�m�G��H����W��_�D��e�w�u�u�w��G��I����V��^�D��d�d�d�d�f�l�G���Y���D��^�E��e�d�e�d�f�m�F��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�e�e�y�]�}�W��I����V��_�D��e�d�d�d�f�l�F��I���F�^�E��e�e�e�e�f�m�F��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�e�u�}�W���[����V��^�D��e�e�e�d�f�l�F��H����FǻN��E��e�e�e�e�f�l�G��H����W��_�E��y�_�u�u�g�m�G��I����W��^�D��d�d�d�d�g�l�[�ԜY���V��^�E��e�e�e�d�f�l�F��H����W�d��U���e�e�e�e�g�m�G��H����W��_�D��d�w�u�u�w��G��I����V��_�E��d�d�d�d�f�l�F���Y���D��^�E��e�d�d�e�g�l�F��H����W��L����u�e�e�e�g�m�G��H����W��_�D��d�e�e�y�]�}�W��I����V��_�D��e�d�d�d�f�l�F��H���F�^�E��e�e�e�e�f�l�G��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�d�u�}�W���[����V��^�D��e�e�e�d�f�l�F��H����FǻN��E��e�e�e�e�f�m�G��I����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�f�m�[�ԜY���V��^�E��d�e�d�e�f�l�F��H����W�d��U���e�e�e�e�g�m�F��I����W��_�D��e�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�F���Y���D��^�E��e�d�e�d�f�m�F��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�d�e�y�]�}�W��I����V��_�E��d�d�d�d�f�l�F��H���F�^�E��e�e�e�d�g�l�G��H����W��_�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�D��d�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�f�m�F��H����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�F��I����V��^�E��d�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�F���Y���D��^�E��e�d�e�e�f�l�G��I����V��L����u�e�e�e�g�m�G��I����W��^�E��e�d�e�y�]�}�W��I����V��_�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�d�g�m�G��I����V��_�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��^�D��d�d�e�e�g�m�G��I����FǻN��E��e�e�e�e�f�l�F��I����V��^�D��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�f�l�[�ԜY���V��^�E��e�d�e�d�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�l�G���Y���D��^�E��e�d�d�e�g�m�G��I����W��L����u�e�e�e�g�m�G��I����W��^�E��e�e�d�y�]�}�W��I����V��_�D��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�f�l�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�d�u�}�W���[����V��^�D��d�d�e�e�g�m�G��H����FǻN��E��e�e�e�e�f�m�G��H����V��^�D��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�f�l�[�ԜY���V��^�E��d�d�d�e�g�m�G��I����W�d��U���e�e�e�e�g�m�F��I����V��^�E��d�w�u�u�w��G��I����V��^�E��e�e�e�e�g�l�F���Y���D��^�E��e�e�d�e�g�m�G��I����W��L����u�e�e�e�g�m�G��I����W��^�E��e�d�d�y�]�}�W��I����V��^�D��d�e�e�e�g�m�F��I���F�^�E��e�e�e�d�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��d�e�d�e�g�m�G��I����FǻN��E��e�e�e�e�g�l�F��H����V��^�E��y�_�u�u�g�m�G��I����W��_�E��e�e�e�d�g�m�[�ԜY���V��^�E��e�d�d�d�g�m�G��I����W�d��U���e�e�e�e�g�m�G��I����V��^�E��d�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�F���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��d�d�e�y�]�}�W��H����W��_�E��d�e�e�e�g�m�F��H���F�_�D��d�d�d�d�g�m�F��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�e�u�}�W���[����W��_�D��d�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��I����V��^�D��y�_�u�u�f�l�F��H����W��^�E��e�e�e�d�f�m�[�ԜY���W��_�D��e�e�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�G��H����V��^�E��d�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�F���Y���D��_�D��d�d�e�d�g�m�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��d�d�d�y�]�}�W��H����W��^�D��d�e�e�e�g�m�F��H���F�_�D��d�d�d�d�g�l�F��I����V��_�W���u�u�w�d�f�l�F��H����V��^�E��e�e�d�e�u�}�W���[����W��_�E��d�e�d�e�g�m�G��H����FǻN��D��d�d�d�d�g�m�G��I����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�d�g�m�[�ԜY���W��_�D��e�e�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�G��H����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�l�G���Y���D��_�D��d�e�e�e�f�m�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��d�d�d�y�]�}�W��H����W��_�E��d�e�e�e�g�m�F��H���F�_�D��d�d�e�d�g�l�G��I����V��_�W���u�u�w�d�f�l�F��I����V��^�E��e�e�e�d�u�}�W���[����W��_�D��d�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��I����V��^�D��y�_�u�u�f�l�F��H����W��_�E��e�e�e�d�f�m�[�ԜY���W��_�D��e�e�d�e�g�m�G��I����V�d��U���d�d�d�d�f�m�G��I����V��^�E��e�w�u�u�w��F��H����V��_�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�g�m�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��d�d�e�y�]�}�W��H����W��^�D��d�e�e�e�g�m�F��I���F�_�D��d�d�e�d�g�l�F��I����V��^�W���u�u�w�d�f�l�F��I����W��^�E��e�e�e�d�u�}�W���[����W��_�E��d�e�e�e�g�m�G��I����FǻN��D��d�d�d�d�g�m�G��H����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�d�g�l�[�ԜY���W��_�D��d�e�d�e�g�m�G��I����V�d��U���d�d�d�d�f�m�G��H����V��^�E��d�w�u�u�w��F��H����V��_�E��e�e�e�e�g�l�F���Y���D��_�D��d�e�d�d�f�m�G��I����W��L����u�d�d�d�f�l�F��H����V��^�E��e�d�d�y�]�}�W��H����W��^�E��d�e�e�e�g�m�G��I���F�_�D��d�d�e�e�f�m�F��I����V��_�W���u�u�w�d�f�l�F��I����W��^�E��e�e�d�d�u�}�W���[����W��_�E��e�e�e�e�g�m�G��H����FǻN��D��d�d�d�d�g�m�F��H����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��e�e�d�d�g�m�G��I����W�d��U���d�d�d�d�f�m�G��I����V��^�E��d�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��e�d�d�d�g�m�G��I����V��L����u�d�d�d�f�l�G��H����W��^�E��e�e�d�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��I���F�_�D��d�d�d�d�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�D��d�d�e�d�f�l�F��H����FǻN��D��d�d�d�e�f�l�F��I����W��_�D��y�_�u�u�f�l�F��H����W��_�D��d�d�d�d�f�m�[�ԜY���W��_�D��e�e�e�e�f�l�F��H����W�d��U���d�d�d�d�f�m�G��I����W��_�D��d�w�u�u�w��F��H����V��^�D��d�d�d�d�f�l�G���Y���D��_�D��d�e�e�d�f�m�F��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�d�e�y�]�}�W��H����W��^�D��d�d�d�d�f�l�F��H���F�_�D��d�d�e�e�f�m�F��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��d�d�e�d�u�}�W���[����W��_�E��d�e�d�d�f�l�F��I����FǻN��D��d�d�d�d�g�l�G��H����W��_�E��y�_�u�u�f�l�F��H����W��_�D��d�d�d�e�f�l�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����V�d��U���d�d�d�d�f�m�F��H����W��_�D��e�w�u�u�w��F��H����V��_�D��d�d�d�d�f�l�F���Y���D��_�D��d�e�d�e�f�l�F��H����W��L����u�d�d�d�f�l�F��H����V��_�D��e�e�d�y�]�}�W��H����W��^�D��e�d�d�d�f�l�G��H���F�_�D��d�d�e�e�g�l�F��H����W��_�W���u�u�w�d�f�l�F��I����W��_�D��d�d�e�e�u�}�W���[����W��_�D��e�d�e�d�f�l�F��I����FǻN��D��d�d�d�d�f�l�G��I����W��_�E��y�_�u�u�f�l�F��H����V��^�D��d�d�d�e�g�l�[�ԜY���W��_�D��d�d�e�d�f�l�F��H����V�d��U���d�d�d�d�f�m�F��I����W��_�E��d�w�u�u�w��F��H����V��_�D��d�d�d�d�g�l�F���Y���D��_�D��d�e�e�e�g�l�F��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�d�e�y�]�}�W��H����W��^�E��d�d�d�d�f�l�F��I���F�_�D��d�d�d�e�f�l�F��H����W��^�W���u�u�w�d�f�l�F��H����V��_�D��d�e�d�e�u�}�W���[����W��_�E��e�e�e�d�f�l�F��I����FǻN��D��d�d�d�d�g�l�F��I����W��^�D��y�_�u�u�f�l�F��H����V��_�D��d�d�d�d�f�l�[�ԜY���W��_�D��e�e�d�d�f�l�F��H����W�d��U���d�d�d�d�f�l�G��I����W��_�E��e�w�u�u�w��F��H����W��_�E��d�d�d�d�g�m�F���Y���D��_�D��d�d�d�d�g�l�F��H����V��L����u�e�e�e�g�m�G��I����V��_�D��d�e�d�y�]�}�W��I����V��^�D��e�d�d�d�f�l�F��I���F�^�E��e�e�e�e�f�m�G��H����W��^�W���u�u�w�e�g�m�G��I����V��_�D��d�e�d�d�u�}�W���[����V��^�E��e�e�e�d�f�l�F��H����FǻN��E��e�e�e�e�g�l�F��I����W��^�D��y�_�u�u�g�m�G��I����V��_�D��d�d�d�e�f�l�[�ԜY���V��^�E��e�e�d�d�f�l�F��H����W�d��U���e�e�e�e�g�m�F��H����W��_�E��e�w�u�u�w��G��I����V��^�E��d�d�d�d�g�l�G���Y���D��^�E��e�d�d�d�f�l�F��H����W��L����u�e�e�e�g�m�G��I����W��_�D��e�d�e�y�]�}�W��I����V��^�E��d�d�d�d�f�l�G��H���F�^�E��e�e�d�d�g�m�F��H����W��^�W���u�u�w�e�g�m�G��H����W��_�D��d�e�d�d�u�}�W���[����V��^�E��d�d�e�d�f�l�F��H����FǻN��E��e�e�e�e�f�m�F��H����W��^�E��y�_�u�u�g�m�G��I����W��_�D��d�d�d�e�g�l�[�ԜY���V��^�E��d�e�d�d�f�l�F��H����W�d��U���e�e�e�e�g�l�F��H����W��_�E��d�w�u�u�w��G��I����V��^�D��d�d�d�d�g�l�G���Y���D��^�E��d�e�e�d�g�m�F��H����W��L����u�e�e�e�g�m�F��H����W��_�D��e�d�e�y�]�}�W��I����V��^�E��d�d�d�d�f�l�G��H���F�^�E��e�e�e�d�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�e�d�d�u�}�W���[����V��^�D��d�d�d�d�f�l�F��H����FǻN��E��e�e�e�d�f�l�G��I����W��^�D��y�_�u�u�g�m�G��I����V��_�D��d�d�d�d�g�m�[�ԜY���V��^�E��d�e�e�d�f�l�F��H����W�d��U���e�e�e�e�g�m�F��I����W��_�E��e�w�u�u�w��G��I����W��_�E��d�d�d�d�g�m�F���Y���D��^�E��d�e�d�e�f�m�F��H����V��L����u�e�e�e�g�m�F��H����V��_�D��d�d�e�y�]�}�W��I����V��^�D��e�d�d�d�f�l�F��I���F�^�E��e�e�d�d�g�l�G��H����W��_�W���u�u�w�e�g�m�G��H����V��_�D��d�e�d�e�u�}�W���[����V��^�D��d�d�e�d�f�l�F��H����FǻN��E��e�e�e�d�f�l�G��I����W��^�E��y�_�u�u�g�m�G��I����W��_�D��d�d�d�d�f�m�[�ԜY���V��^�E��d�e�d�e�f�l�F��H����V�d��U���e�e�e�e�g�l�F��H����W��_�E��d�w�u�u�w��G��I����W��^�E��d�d�d�d�f�m�G���Y���D��^�E��d�d�d�e�f�m�F��H����V��L����u�e�e�e�g�m�G��I����V��_�D��e�d�e�y�]�}�W��I����V��^�E��e�d�d�d�f�l�G��I���F�^�E��e�d�e�e�f�m�G��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�e�u�}�W���[����V��_�E��e�e�e�d�f�l�F��H����FǻN��E��e�e�e�e�g�l�F��I����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�e�f�l�[�ԜY���V��^�D��d�e�e�e�f�l�F��H����W�d��U���e�e�e�e�f�m�F��H����W��_�D��e�w�u�u�w��G��I����V��_�E��d�d�d�d�f�m�F���Y���D��^�E��e�e�e�d�g�m�F��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�e�e�y�]�}�W��I����V��^�D��d�d�d�d�f�l�F��I���F�^�E��e�d�e�d�f�l�F��H����W��_�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��_�E��d�d�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�F��H����V��^�D��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�D��d�e�d�d�g�m�G��I����W�d��U���e�e�e�e�f�m�F��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�d�e�f�l�G��I����V��L����u�e�e�e�g�m�G��H����V��^�E��d�d�d�y�]�}�W��I����V��^�E��d�e�e�e�g�m�F��H���F�^�E��e�d�e�e�f�l�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�e�u�}�W���[����V��^�D��e�d�d�e�g�m�G��H����FǻN��E��e�e�e�d�f�l�G��I����V��_�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�f�m�[�ԜY���V��^�E��d�e�e�e�g�m�G��I����W�d��U���e�e�e�e�g�l�G��H����V��^�D��e�w�u�u�w��G��I����W��_�D��e�e�e�e�f�l�G���Y���D��^�E��d�e�d�d�f�m�G��I����W��L����u�e�e�e�g�m�F��H����W��^�E��d�e�d�y�]�}�W��I����V��^�E��d�e�e�e�g�m�F��H���F�^�E��e�e�d�e�f�m�G��I����V��_�W���u�u�w�e�g�m�G��H����W��^�E��e�d�d�e�u�}�W���[����V��^�D��d�e�d�e�g�m�G��H����FǻN��E��e�e�e�d�f�m�F��I����V��_�D��y�_�u�u�g�m�G��I����W��_�E��e�e�e�d�f�l�[�ԜY���V��^�E��e�d�e�d�g�m�G��H����V�d��U���e�e�e�e�g�m�F��H����V��^�E��e�w�u�u�w��G��I����V��_�E��e�e�e�e�g�m�F���Y���D��^�E��d�e�d�d�f�l�G��I����W��L����u�e�e�e�g�m�F��I����W��^�E��e�e�d�y�]�}�W��I����V��_�E��e�e�e�e�g�l�G��H���F�^�E��e�e�d�e�f�l�G��I����W��_�W���u�u�w�e�g�m�G��H����W��^�E��e�e�e�e�u�}�W���[����V��^�E��d�d�d�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�D��y�_�u�u�g�m�G��I����V��^�E��e�e�d�d�f�l�[�ԜY���V��^�E��d�e�e�e�g�m�G��H����V�d��U���e�e�e�e�g�m�G��I����V��^�E��d�w�u�u�w��G��I����V��^�D��e�e�e�e�g�l�G���Y���D��^�E��e�e�e�d�f�l�G��I����W��L����u�e�e�e�g�m�G��H����V��^�E��d�d�d�y�]�}�W��I����V��^�E��e�e�e�e�g�l�G��I���F�_�D��d�d�d�d�g�l�F��I����W��^�W���u�u�w�d�f�l�F��H����W��^�E��e�d�e�d�u�}�W���[����W��_�E��d�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�g�l�F��I����V��_�D��y�_�u�u�f�l�F��H����V��_�E��e�e�d�e�f�l�[�ԜY���W��_�D��d�d�d�e�g�m�G��H����V�d��U���d�d�d�d�f�m�G��I����V��^�D��d�w�u�u�w��F��H����V��^�E��e�e�e�e�f�l�G���Y���D��_�D��d�e�d�d�g�m�G��I����W��L����u�d�d�d�f�l�F��I����W��^�E��e�e�d�y�]�}�W��H����W��_�D��e�e�e�e�g�l�G��H���F�_�D��d�d�d�e�f�m�F��I����W��^�W���u�u�w�d�f�l�F��H����W��^�E��e�d�d�e�u�}�W���[����W��_�E��e�d�d�e�g�m�G��H����FǻN��D��d�d�d�e�f�l�F��H����V��_�E��y�_�u�u�f�l�F��H����V��^�E��e�e�d�e�g�l�[�ԜY���W��_�D��e�d�d�d�g�m�G��H����W�d��U���d�d�d�d�f�m�F��I����V��^�D��e�w�u�u�w��F��H����V��^�E��e�e�e�e�f�m�F���Y���D��_�D��d�d�d�d�f�m�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�d�e�y�]�}�W��H����W��_�D��e�e�e�e�g�l�G��H���F�_�D��d�e�d�d�g�m�G��I����W��_�W���u�u�w�d�f�l�F��H����V��^�E��e�d�e�d�u�}�W���[����W��^�E��e�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��I����V��_�E��y�_�u�u�f�l�F��H����W��^�E��e�e�d�d�f�l�[�ԜY���W��_�E��d�d�e�e�g�m�G��H����W�d��U���d�d�d�d�g�m�F��H����V��^�E��d�w�u�u�w��F��H����V��_�E��e�e�e�e�g�l�G���Y���D��_�D��e�d�d�d�g�l�G��I����V��L����u�d�d�d�f�l�G��I����V��^�E��d�d�d�y�]�}�W��H����W��_�D��e�e�e�e�g�l�F��H���F�_�D��d�e�d�d�f�m�G��I����W��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�d�d�u�}�W���[����W��^�E��e�d�d�e�g�m�G��H����FǻN��D��d�d�d�e�f�l�F��H����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�d�e�f�m�[�ԜY���W��_�E��e�d�e�d�g�m�G��H����W�d��U���d�d�d�d�g�m�G��I����V��^�E��e�w�u�u�w��F��H����V��_�E��e�e�e�e�f�l�G���Y���D��_�D��e�e�e�d�f�l�G��I����W��L����u�d�d�d�f�l�G��I����W��^�E��d�d�e�y�]�}�W��H����W��^�E��d�e�e�e�g�m�F��H���F�_�D��d�e�e�e�f�m�F��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�d�d�e�u�}�W���[����W��_�D��d�e�d�e�g�m�G��H����FǻN��D��d�d�e�d�f�m�G��H����V��_�D��y�_�u�u�f�l�F��I����V��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��e�d�e�d�g�m�G��I����V�d��U���d�d�d�d�f�l�G��H����V��^�E��e�w�u�u�w��F��H����W��^�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�d�f�l�G��I����V��L����u�d�d�d�f�m�F��I����W��^�E��e�d�e�y�]�}�W��H����V��_�D��e�e�e�e�g�m�G��H���F�_�D��d�d�d�e�f�m�G��I����V��^�W���u�u�w�d�f�l�F��H����V��_�D��d�d�d�d�u�}�W���[����W��_�D��e�e�e�d�f�l�F��H����FǻN��D��d�d�e�d�f�m�F��H����W��_�D��y�_�u�u�f�l�F��I����W��^�D��d�d�d�d�g�l�[�ԜY���W��_�D��e�e�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�G��H����W��_�D��d�w�u�u�w��F��H����W��^�D��d�d�d�d�f�m�F���Y���D��_�D��d�d�e�e�f�m�F��H����W��L����u�d�d�d�f�m�F��H����W��_�D��d�e�d�y�]�}�W��H����W��^�E��e�d�d�d�f�l�F��H���F�_�D��d�e�e�e�f�m�G��H����W��^�W���u�u�w�d�f�l�F��I����V��_�D��d�e�d�d�u�}�W���[����W��^�E��d�d�d�d�f�l�F��I����FǻN��D��d�d�d�e�g�l�F��I����W��^�E��y�_�u�u�f�l�F��H����V��^�D��d�d�e�d�f�l�[�ԜY���W��_�E��e�d�d�d�f�l�F��I����V�d��U���d�d�d�d�g�m�F��I����W��_�D��d�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�F���Y���D��_�D��e�e�d�d�f�l�F��H����W��L����u�d�d�d�f�l�G��I����V��_�D��e�d�d�y�]�}�W��H����W��_�E��e�d�d�d�f�m�G��I���F�_�D��d�e�d�e�f�l�G��H����V��_�W���u�u�w�d�f�l�F��H����V��_�D��d�e�e�d�u�}�W���[����W��^�E��d�e�d�d�f�l�F��I����FǻN��D��d�d�d�d�g�l�G��H����W��^�D��y�_�u�u�f�l�F��H����V��^�D��d�d�e�e�g�m�[�ԜY���W��_�E��d�d�e�e�f�l�F��I����V�d��U���d�d�d�d�g�l�G��I����W��_�E��d�w�u�u�w��F��H����W��_�D��d�d�d�e�f�l�G���Y���D��_�D��d�d�e�d�f�l�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�e�y�]�}�W��H����W��^�E��e�d�d�d�f�l�F��I���F�_�D��d�d�e�d�f�m�F��H����W��_�W���u�u�w�d�f�l�F��I����W��_�D��e�d�d�d�u�}�W���[����W��_�E��d�d�e�d�f�l�G��I����FǻN��D��d�d�d�e�g�m�F��I����W��_�D��y�_�u�u�f�l�F��H����W��^�D��d�d�d�e�g�m�[�ԜY���W��_�D��d�d�e�e�f�l�F��H����W�d��U���d�d�d�d�f�m�F��H����W��_�E��d�w�u�u�w��F��H����V��^�D��d�d�d�e�g�m�F���Y���D��_�D��d�d�d�e�f�l�F��H����V��L����u�d�d�d�f�l�F��I����W��_�D��d�e�e�y�]�}�W��H����W��_�E��e�d�d�d�f�l�F��I���F�^�E��e�e�e�e�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��e�e�d�d�u�}�W���[����V��^�D��e�e�d�d�f�l�G��H����FǻN��E��e�e�e�e�g�m�G��I����W��^�E��y�_�u�u�g�m�G��I����W��_�D��d�d�d�e�f�m�[�ԜY���V��^�E��d�e�d�e�f�l�F��H����W�d��U���e�e�e�e�g�m�G��I����W��_�E��d�w�u�u�w��G��I����V��^�E��d�d�d�e�g�m�F���Y���D��^�E��d�d�d�d�g�m�F��H����V��L����u�e�e�e�g�m�F��I����W��_�D��e�e�d�y�]�}�W��I����V��_�E��e�d�d�d�f�l�G��I���F�^�E��e�d�e�e�g�m�G��H����W��^�W���u�u�w�e�g�m�G��I����V��_�D��e�e�e�e�u�}�W���[����V��_�D��d�e�d�d�f�l�G��I����FǻN��E��e�e�e�e�g�l�F��I����W��^�E��y�_�u�u�g�m�G��I����V��_�D��d�d�d�e�g�l�[�ԜY���V��^�D��d�e�d�e�f�l�F��H����V�d��U���e�e�e�e�f�m�F��H����W��_�E��d�w�u�u�w��G��I����V��^�D��d�d�d�e�g�m�G���Y���D��^�E��d�e�e�e�g�m�F��H����V��L����u�e�e�e�g�m�F��I����W��_�D��e�d�d�y�]�}�W��I����V��_�D��d�d�d�d�f�l�G��I���F�^�E��e�e�e�e�f�l�G��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��e�e�d�e�u�}�W���[����V��^�D��e�d�d�d�f�l�G��H����FǻN��E��e�e�d�e�g�m�F��H����W��^�E��y�_�u�u�g�m�G��H����W��_�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�e�d�d�f�l�F��H����V�d��U���e�e�e�e�g�m�G��I����W��_�E��d�w�u�u�w��G��I����V��^�D��d�d�d�e�g�l�F���Y���D��^�E��d�d�d�d�f�m�F��H����V��L����u�e�e�e�g�l�F��I����V��_�D��e�d�e�y�]�}�W��I����W��^�D��e�d�d�d�f�l�G��I���F�^�E��e�e�d�e�f�m�F��H����W��_�W���u�u�w�e�g�m�G��H����V��_�D��e�d�e�d�u�}�W���[����V��_�E��e�d�e�d�f�l�G��I����FǻN��E��e�e�d�e�g�l�F��I����W��_�D��y�_�u�u�g�m�G��H����W��_�D��d�d�e�e�g�l�[�ԜY���V��^�D��d�e�d�e�f�l�F��I����W�d��U���e�e�e�e�f�l�G��H����W��_�E��e�w�u�u�w��G��I����W��_�E��d�d�d�d�g�m�F���Y���D��^�E��e�d�e�d�g�l�F��H����V��L����u�e�e�e�g�l�G��H����V��_�D��d�d�d�y�]�}�W��I����W��_�E��d�d�d�d�f�m�G��I���F�^�E��e�d�e�e�f�l�G��H����V��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�e�e�u�}�W���[����V��_�E��e�e�d�d�f�l�F��I����FǻN��E��e�e�d�d�f�m�G��I����W��_�D��y�_�u�u�g�m�G��H����V��_�D��d�d�d�e�f�l�[�ԜY���V��^�D��e�d�e�d�f�l�F��H����V�d��U���e�e�e�e�f�m�F��I����W��_�E��d�w�u�u�w��G��I����V��^�D��d�d�d�d�g�l�F���Y���D��^�E��d�d�d�e�f�l�F��H����V��L����u�e�e�e�g�l�F��H����V��_�D��e�e�d�y�]�}�W��I����W��^�E��d�d�d�d�f�l�F��H���F�^�E��e�d�d�e�g�m�F��H����W��^�W���u�u�w�e�g�m�G��H����V��^�E��e�e�e�e�u�}�W���[����V��_�E��e�e�e�e�g�m�G��H����FǻN��E��e�e�d�d�f�l�F��I����V��^�E��y�_�u�u�g�m�G��H����W��^�E��e�e�e�d�g�m�[�ԜY���V��^�D��d�e�e�e�g�m�G��I����V�d��U���e�e�e�e�f�m�F��H����V��^�D��e�w�u�u�w��G��I����V��_�E��e�e�e�e�f�m�G���Y���D��^�E��d�d�e�e�f�l�G��I����W��L����u�e�e�e�g�l�F��H����V��^�E��e�e�d�y�]�}�W��I����W��^�D��e�e�e�e�g�l�G��I���F�^�E��e�d�e�e�g�m�F��I����W��^�W���u�u�w�e�g�m�G��H����V��^�E��e�e�d�d�u�}�W���[����V��_�D��d�d�d�e�g�m�G��I����FǻN��E��e�e�d�e�f�m�G��I����V��_�E��y�_�u�u�g�m�G��H����V��_�E��e�e�d�d�g�l�[�ԜY���V��^�D��e�d�d�d�g�m�G��H����V�d��U���e�e�e�e�f�m�F��I����V��^�E��e�w�u�u�w��G��I����V��_�E��e�e�e�d�g�l�G���Y���D��^�E��e�e�e�d�f�l�G��I����V��L����u�e�e�e�g�l�F��H����W��^�E��d�d�e�y�]�}�W��I����W��_�E��d�e�e�e�g�m�G��I���F�^�E��e�e�d�d�f�l�F��I����V��_�W���u�u�w�e�g�m�G��I����V��^�E��d�d�e�e�u�}�W���[����V��^�D��d�d�e�e�g�m�F��H����FǻN��E��e�e�d�d�g�l�F��I����V��^�E��y�_�u�u�g�m�G��H����V��_�E��e�e�d�e�g�l�[�ԜY���V��^�E��d�e�d�e�g�m�G��H����V�d��U���e�e�e�e�g�l�G��I����V��^�E��e�w�u�u�w��G��I����V��_�E��e�e�e�d�f�m�G���Y���D��^�E��e�e�e�d�f�m�G��I����V��L����u�e�e�e�g�m�F��H����V��^�E��e�d�e�y�]�}�W��I����V��^�E��d�e�e�e�g�l�F��I���F�^�E��e�d�e�e�f�m�G��I����W��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�e�u�}�W���[����V��_�D��d�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�l�G��I����V��^�D��y�_�u�u�g�m�G��I����V��^�E��e�d�e�d�g�m�[�ԜY���V��^�D��e�d�e�d�g�m�G��I����W�d��U���e�e�e�e�g�l�G��I����V��_�E��e�w�u�u�w��G��I����V��_�D��e�e�e�e�f�m�G���Y���D��^�E��d�e�e�d�f�l�G��I����V��L����u�e�e�e�g�m�G��I����W��^�D��e�e�e�y�]�}�W��I����V��^�D��d�e�e�e�f�m�G��I���F�^�E��e�e�e�e�f�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�d�e�e�u�}�W���[����W��_�E��e�d�d�e�g�m�G��H����FǻN��D��d�d�d�d�f�m�G��I����V��_�D��y�_�u�u�f�l�F��H����W��_�E��e�d�e�d�f�m�[�ԜY���W��_�D��e�e�d�e�g�m�G��H����W�d��U���d�d�d�d�f�m�F��H����V��_�E��d�w�u�u�w��F��H����V��^�D��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�e�g�m�G��I����V��L����u�d�d�d�f�l�F��H����V��^�D��e�d�d�y�]�}�W��H����W��^�D��d�e�e�e�f�l�G��I���F�_�D��d�e�d�e�f�l�F��I����W��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�d�e�u�}�W���[����W��^�E��d�e�e�e�g�m�G��H����FǻN��D��d�d�e�d�f�m�F��H����V��^�D��y�_�u�u�f�l�F��I����W��_�E��e�d�d�e�f�m�[�ԜY���W��_�D��e�e�d�e�g�m�G��H����W�d��U���d�d�d�d�f�l�F��I����V��_�E��d�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��e�d�d�e�f�m�G��I����W��L����u�d�d�d�f�m�G��I����V��^�D��d�d�e�y�]�}�W��H����V��^�E��d�e�e�e�f�m�F��H���F�_�D��d�e�e�d�g�l�G��I����V��_�W���u�u�w�d�f�l�F��I����V��^�E��e�d�e�d�u�}�W���[����W��^�D��d�e�e�e�g�m�G��H����FǻN��D��d�d�e�e�g�m�G��H����V��_�E��y�_�u�u�f�l�F��I����W��^�E��e�d�e�e�f�l�[�ԜY���W��_�D��d�e�d�d�g�m�G��I����V�d��U���d�d�d�e�f�l�F��I����V��_�E��d�w�u�u�w��F��H����V��^�D��e�e�e�e�g�m�G���Y���D��_�D��d�e�e�e�f�m�G��I����W��L����u�d�d�d�f�l�G��I����V��^�D��e�e�e�y�]�}�W��H����W��^�E��d�e�e�e�f�m�G��H���F�_�D��e�d�e�d�g�l�G��I����W��^�W���u�u�w�d�f�l�G��I����W��^�E��d�d�e�d�u�}�W���[����W��^�D��d�e�e�e�g�m�F��H����FǻN��D��d�d�d�d�g�l�G��H����V��_�E��y�_�u�u�f�l�F��H����W��_�E��e�e�d�d�g�l�[�ԜY���W��_�E��e�d�e�e�g�m�G��H����W�d��U���d�d�d�e�g�m�G��H����V��^�E��d�w�u�u�w��F��H����W��^�D��e�e�e�d�f�l�F���Y���D��_�D��e�e�d�e�g�l�G��I����V��L����u�d�d�d�f�l�G��H����W��^�E��e�e�e�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��I���F�_�D��e�e�e�e�g�l�F��I����V��_�W���u�u�w�d�f�l�G��I����V��^�E��d�e�d�d�u�}�W���[����W��^�E��e�e�d�e�g�m�F��I����FǻN��D��d�d�e�d�f�m�G��I����V��_�D��y�_�u�u�f�l�F��I����V��_�E��e�e�d�e�g�l�[�ԜY���W��_�D��d�e�e�d�g�m�G��H����W�d��U���d�d�d�e�f�l�G��I����V��^�E��e�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�d�d�f�l�G��I����W��L����u�d�d�d�f�m�F��H����W��^�E��e�d�e�y�]�}�W��H����V��_�D��e�e�e�e�g�m�G��I���F�_�D��e�d�e�d�g�l�G��I����V��^�W���u�u�w�d�f�l�G��I����V��^�E��e�e�e�d�u�}�W���[����W��_�D��d�e�d�d�f�l�F��H����FǻN��D��d�d�e�d�f�m�G��H����W��_�E��y�_�u�u�f�l�F��I����W��^�D��d�d�d�d�f�m�[�ԜY���W��_�D��e�e�e�e�f�l�F��H����W�d��U���d�d�d�e�f�l�G��H����W��_�E��d�w�u�u�w��F��H����W��^�E��d�d�d�d�f�m�G���Y���D��_�D��d�e�d�e�g�m�F��H����W��L����u�d�d�d�f�m�F��H����V��_�D��d�e�e�y�]�}�W��H����V��_�D��d�d�d�d�f�m�G��I���F�_�D��e�e�e�e�f�l�F��H����W��_�W���u�u�w�d�f�l�G��I����W��_�D��e�d�e�e�u�}�W���[����W��^�D��e�d�d�d�f�l�G��I����FǻN��D��d�d�d�e�g�m�F��I����W��^�D��y�_�u�u�f�l�F��H����W��^�D��d�d�d�e�g�m�[�ԜY���W��_�E��d�e�e�e�f�l�F��I����V�d��U���d�d�d�e�g�m�G��I����W��_�D��e�w�u�u�w��F��H����V��^�D��d�d�d�e�g�l�F���Y���D��_�D��d�e�e�d�g�m�F��H����V��L����u�d�d�d�f�l�F��I����W��_�D��e�d�d�y�]�}�W��H����W��^�D��e�d�d�d�g�l�F��I���F�_�D��e�d�e�e�g�l�F��H����W��^�W���u�u�w�d�f�l�G��H����W��_�D��d�e�d�d�u�}�W���[����W��_�D��d�d�e�d�f�l�F��I����FǻN��D��d�d�d�d�g�l�F��H����W��^�D��y�_�u�u�f�l�F��H����V��_�D��d�e�e�d�g�l�[�ԜY���W��_�D��e�d�e�d�f�l�F��I����W�d��U���d�d�d�d�g�m�F��I����W��^�D��e�w�u�u�w��F��H����W��_�E��d�d�d�d�g�m�G���Y���D��_�D��e�d�e�d�g�l�F��H����W��L����u�d�d�d�f�m�F��I����V��_�E��d�d�d�y�]�}�W��H����V��^�D��d�d�d�d�g�l�F��I���F�_�D��d�d�e�e�g�m�G��H����W��^�W���u�u�w�d�f�l�F��I����V��_�D��e�d�e�e�u�}�W���[����W��_�D��d�d�e�d�f�l�G��I����FǻN��D��d�d�e�d�f�l�F��H����W��^�D��y�_�u�u�f�l�F��I����V��_�D��d�e�d�e�f�m�[�ԜY���W��_�E��d�e�e�d�f�l�F��I����W�d��U���d�d�d�d�g�l�F��H����W��^�D��d�w�u�u�w��F��H����V��_�D��d�d�d�e�f�l�F���Y���D��_�D��d�e�d�d�g�m�F��H����V��L����u�d�d�d�f�l�G��I����V��_�E��d�d�e�y�]�}�W��H����W��^�E��d�d�d�d�g�m�F��I���F�_�D��d�d�e�e�g�l�F��H����V��^�W���u�u�w�d�f�l�F��H����V��_�D��e�e�d�d�u�}�W���[����V��^�E��e�e�e�d�f�l�G��I����FǻN��E��e�e�e�e�g�m�G��I����W��^�E��y�_�u�u�g�m�G��I����V��_�D��d�d�d�d�g�l�[�ԜY���V��^�E��e�e�d�e�f�l�F��H����V�d��U���e�e�e�e�f�m�G��H����W��_�D��e�w�u�u�w��G��I����W��_�D��d�d�e�d�f�m�G���Y���D��^�E��d�e�e�d�g�m�F��I����W��L����u�e�e�e�g�m�F��H����W��_�D��e�d�d�y�]�}�W��I����W��^�E��d�d�d�d�f�l�G��I���F�^�E��e�e�d�e�f�m�G��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�d�u�}�W���[����V��^�E��d�d�d�d�f�m�F��H����FǻN��E��e�e�d�e�g�m�F��H����V��_�D��y�_�u�u�g�m�G��H����W��^�D��d�d�d�e�f�m�[�ԜY���V��^�D��d�e�e�d�f�l�F��H����V�d��U���e�e�e�e�f�l�F��I����W��_�D��d�w�u�u�w��G��I����V��_�D��d�d�e�d�f�m�G���Y���D��^�E��e�e�d�d�g�l�F��I����W��L����u�e�e�e�g�m�F��H����W��_�D��d�d�d�y�]�}�W��I����V��^�D��d�d�d�d�g�m�G��I���F�^�E��d�d�e�d�f�l�F��H����V��^�W���u�u�w�e�g�m�F��H����W��_�D��e�e�d�d�u�}�W���[����V��_�E��e�e�e�d�f�l�G��I����FǻN��E��e�e�e�d�g�m�G��H����W��^�E��y�_�u�u�g�m�G��H����V��_�D��d�e�e�e�g�l�[�ԜY���V��^�E��e�d�e�e�f�l�F��I����W�d��U���e�e�e�d�g�m�G��H����W��^�D��e�w�u�u�w��G��I����V��_�E��d�d�d�e�f�l�G���Y���D��^�E��d�d�e�e�g�m�F��H����V��L����u�e�e�e�g�l�G��H����V��_�E��d�e�d�y�]�}�W��I����W��^�D��e�d�d�d�g�l�F��I���F�^�E��d�d�e�d�g�m�G��H����W��^�W���u�u�w�e�g�m�F��H����V��_�D��e�d�e�e�u�}�W���[����V��_�D��e�e�d�d�f�l�F��I����FǻN��E��e�d�e�e�f�m�F��I����W��^�D��y�_�u�u�g�m�G��I����W��^�D��d�e�e�d�g�l�[�ԜY���V��_�E��d�e�e�e�f�l�F��I����W�d��U���e�e�e�e�g�m�G��H����W��^�D��d�w�u�u�w��G��I����W��^�E��d�d�d�d�g�m�F���Y���D��^�D��d�d�d�d�f�l�F��H����V��L����u�e�e�e�f�m�G��I����V��_�E��e�d�d�y�]�}�W��I����V��_�D��d�d�d�d�g�l�F��I���F�^�E��e�d�d�d�g�l�G��H����V��_�W���u�u�w�e�g�m�G��H����V��_�D��e�e�e�d�u�}�W���[����V��_�E��d�d�e�d�f�l�G��H����FǻN��E��e�d�e�d�f�m�G��H����W��_�E��y�_�u�u�g�m�G��I����W��_�D��d�d�d�e�f�l�[�ԜY���V��_�D��e�d�e�e�f�l�F��H����V�d��U���e�e�e�e�f�l�G��I����W��_�D��d�w�u�u�w��G��I����W��_�D��d�d�d�d�g�m�F���Y���D��^�D��d�d�d�e�g�m�F��H����W��L����u�e�e�e�f�l�G��I����W��_�D��e�d�d�y�]�}�W��I����W��^�D��d�d�d�d�f�l�G��H���F�^�E��e�e�e�d�g�l�F��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�d�d�d�u�}�W���[����V��^�E��d�d�e�d�f�l�F��H����FǻN��E��e�d�d�e�g�m�G��I����V��^�D��y�_�u�u�g�m�G��H����W��_�E��e�e�e�e�g�l�[�ԜY���V��_�E��e�d�d�e�g�m�G��I����V�d��U���e�e�e�e�f�l�F��I����V��^�E��e�w�u�u�w��G��I����W��_�D��e�e�e�e�f�l�G���Y���D��^�D��d�e�d�d�f�l�G��I����W��L����u�e�e�e�f�m�F��H����V��^�E��d�d�d�y�]�}�W��I����V��_�D��d�e�e�e�g�m�G��I���F�^�E��e�d�e�d�f�l�F��I����W��^�W���u�u�w�e�g�m�G��I����W��^�E��d�e�e�d�u�}�W���[����V��_�D��d�d�e�e�g�m�F��H����FǻN��E��e�d�e�e�g�m�F��H����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�d�e�d�f�l�[�ԜY���V��_�E��d�d�d�e�g�m�G��I����V�d��U���e�e�e�e�g�l�F��I����V��_�E��d�w�u�u�w��G��I����V��_�E��e�e�e�e�g�m�F���Y���D��^�D��e�d�d�d�f�m�G��I����W��L����u�e�e�e�f�m�G��H����W��^�D��e�e�d�y�]�}�W��I����V��^�E��e�e�e�e�f�m�F��I���F�^�E��d�d�d�e�f�m�F��I����V��^�W���u�u�w�e�g�m�F��I����V��^�E��d�d�d�d�u�}�W���[����V��_�D��e�e�d�e�g�m�F��I����FǻN��E��e�e�d�e�f�m�F��H����V��_�D��y�_�u�u�g�m�G��H����W��^�E��e�d�d�d�g�l�[�ԜY���V��^�E��d�d�e�d�g�m�G��I����V�d��U���e�e�e�d�g�l�F��H����V��^�E��d�w�u�u�w��G��I����V��_�D��e�e�d�e�f�m�G���Y���D��^�E��d�d�e�e�f�m�G��H����V��L����u�e�e�e�g�m�F��H����V��^�E��d�d�e�y�]�}�W��I����V��^�D��d�e�e�e�g�l�G��H���F�^�E��d�e�d�d�f�m�G��I����W��_�W���u�u�w�e�g�m�F��I����V��^�E��d�e�e�d�u�}�W���[����V��^�E��d�e�d�e�g�l�F��I����FǻN��E��e�e�e�e�g�m�F��H����W��_�D��y�_�u�u�g�m�G��H����V��_�E��e�e�e�d�g�m�[�ԜY���V��^�D��d�e�e�e�g�m�G��H����V�d��U���e�e�e�e�g�l�F��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�d�d�g�l�F���Y���D��^�E��e�e�e�d�g�m�G��H����V��L����u�e�e�e�g�m�F��H����V��^�E��d�e�d�y�]�}�W��I����V��^�E��d�e�e�e�g�l�F��I���F�^�E��e�d�e�e�g�m�G��I����V��_�W���u�u�w�e�g�m�G��H����V��^�E��e�e�d�d�u�}�W���[����V��^�D��d�d�d�e�g�l�G��I����FǻN��E��e�e�e�e�g�m�G��I����W��^�D��y�_�u�u�f�l�F��H����W��^�E��e�d�e�e�f�m�[�ԜY���W��_�D��d�d�d�e�g�m�G��I����V�d��U���d�d�d�d�g�l�G��H����V��_�D��d�w�u�u�w��F��H����W��^�D��e�e�d�e�f�m�F���Y���D��_�D��e�e�e�e�g�m�G��H����W��L����u�d�d�d�f�m�F��H����W��^�D��d�d�e�y�]�}�W��H����V��_�E��e�e�e�e�f�l�G��I���F�_�D��d�e�d�e�g�l�F��I����W��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�d�u�}�W���[����W��_�D��e�d�d�e�g�l�G��I����FǻN��D��d�d�d�d�g�m�G��I����W��^�E��y�_�u�u�f�l�F��H����W��^�E��e�d�e�d�f�l�[�ԜY���W��_�E��e�e�d�d�g�m�G��I����V�d��U���d�d�d�e�g�l�F��I����V��_�D��e�w�u�u�w��F��H����W��^�D��e�e�d�e�f�m�G���Y���D��_�D��d�e�d�d�g�m�G��H����W��L����u�d�d�d�f�m�G��H����V��^�D��e�e�e�y�]�}�W��H����V��^�D��d�e�e�e�f�m�G��H���F�_�D��e�e�d�e�g�l�F��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�e�u�}�W���[����W��_�E��d�d�d�e�g�l�G��I����FǻN��D��d�e�d�e�f�l�F��H����W��_�D��y�_�u�u�f�l�F��H����V��^�E��e�e�d�d�g�m�[�ԜY���W��^�E��e�d�e�d�g�m�G��H����V�d��U���d�d�d�d�g�m�G��I����V��^�E��d�w�u�u�w��F��H����W��^�D��e�e�d�d�g�l�G���Y���D��_�E��e�d�d�e�f�l�G��H����W��L����u�d�d�d�g�m�G��I����W��^�E��e�e�e�y�]�}�W��H����V��^�E��d�e�e�e�g�m�F��H���F�_�D��d�e�e�e�g�m�F��I����V��^�W���u�u�w�d�f�l�F��I����W��^�E��e�d�e�d�u�}�W���[����W��_�D��e�e�d�e�g�l�G��I����FǻN��D��d�e�d�d�g�l�F��I����W��^�D��y�_�u�u�f�l�F��H����V��^�E��e�e�e�d�g�m�[�ԜY���W��^�D��e�d�d�d�g�m�G��I����W�d��U���d�d�d�e�g�l�G��H����V��^�E��d�w�u�u�w��F��H����V��_�D��e�e�e�d�f�l�G���Y���D��_�E��e�e�e�d�g�l�G��I����V��L����u�d�d�d�g�l�G��H����W��^�D��e�e�e�y�]�}�W��H����V��_�E��d�e�e�e�f�m�F��I���F�_�D��e�d�e�d�g�m�G��I����V��_�W���u�u�w�d�f�l�G��I����W��^�E��e�d�d�e�u�}�W���[����W��_�E��e�e�e�e�g�m�G��I����FǻN��D��d�e�e�e�f�l�G��I����V��^�D��y�_�u�u�f�l�F��I����V��^�E��e�d�e�e�g�m�[�ԜY���W��^�E��e�d�d�d�g�m�G��I����W�d��U���d�d�d�e�g�l�G��H����V��^�D��e�w�u�u�w��F��H����V��_�D��e�e�e�d�g�m�F���Y���D��_�E��d�e�e�d�g�m�G��I����V��L����u�d�d�d�g�m�F��I����W��^�E��d�d�d�y�]�}�W��H����V��_�D��d�e�e�e�g�l�F��I���F�_�D��e�e�d�e�g�l�F��I����W��^�W���u�u�w�d�f�l�G��H����V��^�E��e�d�d�e�u�}�W���[����W��^�E��d�e�e�e�g�m�G��H����FǻN��D��d�e�e�e�g�l�F��H����W��_�E��y�_�u�u�f�l�F��I����V��_�D��d�d�d�d�g�l�[�ԜY���W��^�E��e�d�d�d�f�l�F��I����V�d��U���d�d�d�e�g�l�F��I����W��_�E��d�w�u�u�w��F��H����V��_�E��d�d�d�e�f�m�F���Y���D��_�E��d�d�e�e�g�l�F��H����V��L����u�d�d�d�g�m�F��H����W��_�D��d�d�e�y�]�}�W��H����V��^�E��e�d�d�d�f�m�F��I���F�_�D��e�e�d�d�g�m�F��H����W��^�W���u�u�w�d�f�l�G��I����V��_�D��d�e�e�e�u�}�W���[����W��_�E��d�d�d�d�f�l�F��H����FǻN��D��d�e�e�e�f�l�G��I����W��^�D��y�_�u�u�f�l�F��I����W��_�D��d�e�d�e�f�m�[�ԜY���W��^�D��e�e�e�d�f�l�F��H����W�d��U���d�d�d�e�g�m�F��H����W��^�D��d�w�u�u�w��F��H����W��^�D��d�d�d�e�g�l�G���Y���D��_�E��d�e�d�d�f�l�F��I����W��L����u�d�d�d�g�l�F��I����W��_�D��e�e�e�y�]�}�W��H����W��_�E��d�d�d�d�f�m�G��I���F�_�D��e�d�d�d�f�l�F��H����V��^�W���u�u�w�d�f�l�G��H����V��_�D��e�d�d�e�u�}�W���[����W��^�D��e�e�e�d�f�m�G��H����FǻN��D��d�e�e�d�g�m�F��I����V��_�D��y�_�u�u�f�l�F��I����V��_�D��d�d�e�e�f�m�[�ԜY���W��^�D��e�e�d�d�f�l�F��H����W�d��U���d�d�d�d�f�m�G��H����W��^�E��e�w�u�u�w��F��H����V��^�E��d�d�e�d�f�l�G���Y���D��_�E��e�d�d�d�f�m�F��I����W��L����u�d�d�d�g�l�F��H����W��_�E��e�e�d�y�]�}�W��H����W��_�E��d�d�d�d�g�l�G��H���F�_�D��d�d�d�d�g�m�G��H����W��_�W���u�u�w�d�f�l�G��H����W��_�D��e�d�e�e�u�}�W���[����W��^�E��d�e�d�d�f�m�G��H����FǻN��D��d�d�e�e�g�l�G��I����V��^�D��y�_�u�u�f�l�F��I����W��_�D��e�d�d�e�f�m�[�ԜY���W��_�E��d�d�e�e�f�l�G��H����W�d��U���d�d�d�e�g�l�F��I����W��_�E��e�w�u�u�w��F��H����W��_�E��d�d�d�d�f�m�G���Y���D��_�D��d�d�e�d�f�m�F��H����W��L����u�d�d�d�f�m�F��I����V��_�D��e�d�e�y�]�}�W��H����V��^�E��e�d�d�e�f�l�F��H���F�_�D��d�d�e�e�f�m�F��H����W��^�W���u�u�w�d�f�l�F��I����V��_�D��e�e�d�e�u�}�W���[����W��^�E��d�e�e�d�f�l�G��H����FǻN��D��d�d�d�e�f�m�F��I����W��^�E��y�_�u�u�g�m�G��I����V��^�D��e�d�e�d�f�m�[�ԜY���V��^�E��d�e�e�e�f�l�G��I����V�d��U���e�e�e�e�f�m�F��I����W��_�D��d�w�u�u�w��G��I����W��^�D��d�d�d�e�g�l�F���Y���D��^�E��e�d�e�e�g�m�F��H����V��L����u�e�e�e�g�l�G��H����V��_�D��e�d�e�y�]�}�W��I����W��_�D��d�d�d�e�f�m�G��I���F�^�E��d�e�d�e�f�m�F��H����V��_�W���u�u�w�e�g�m�F��H����W��_�D��e�e�e�e�u�}�W���[����V��_�E��d�e�d�d�f�l�G��I����FǻN��E��e�e�d�e�f�l�F��I����W��^�D��y�_�u�u�g�m�G��H����W��_�D��e�d�e�e�f�l�[�ԜY���V��^�D��e�e�e�d�f�l�G��I����W�d��U���e�e�e�e�g�m�G��I����W��_�E��d�w�u�u�w��G��I����V��^�D��d�d�d�e�g�m�G���Y���D��^�D��e�e�e�e�g�m�F��H����W��L����u�e�e�e�f�m�F��H����W��_�D��e�d�d�y�]�}�W��I����W��_�D��e�d�d�e�f�m�G��H���F�^�E��e�d�e�e�f�m�F��H����V��^�W���u�u�w�e�g�m�G��I����W��_�D��e�e�e�d�u�}�W���[����V��^�D��d�d�e�d�f�l�G��I����FǻN��E��e�d�e�d�g�l�F��I����W��_�D��y�_�u�u�g�m�G��I����W��_�D��e�d�d�d�f�l�[�ԜY���V��_�D��e�d�e�d�f�l�G��I����W�d��U���e�e�e�d�g�l�F��H����W��_�E��d�w�u�u�w��G��I����V��_�D��d�d�d�d�f�l�F���Y���D��^�D��d�e�d�e�g�l�F��H����V��L����u�e�e�e�g�m�G��I����V��_�D��d�e�d�y�]�}�W��I����V��^�E��e�d�d�e�f�l�F��H���F�^�E��e�d�e�d�g�m�G��H����V��_�W���u�u�w�e�g�l�G��I����W��_�D��e�d�d�e�u�}�W���[����W��^�E��e�d�d�d�f�m�G��I����FǻN��E��e�e�d�e�f�l�G��I����V��_�E��y�_�u�u�g�m�G��H����W��_�D��d�e�d�d�f�l�[�ԜY���V��^�D��d�d�e�d�f�l�F��I����W�d��U���e�e�d�e�f�m�F��I����W��^�D��d�w�u�u�w��G��H����V��^�D��d�d�e�d�f�m�G���Y���D��^�E��d�e�e�e�g�l�F��I����V��L����u�e�e�e�g�m�F��H����W��_�D��e�e�e�y�]�}�W��I����V��_�E��e�d�d�d�f�l�G��H���F�^�E��d�d�e�e�g�l�G��H����W��^�W���u�u�w�e�g�l�F��H����W��_�D��d�e�d�d�u�}�W���[����W��^�E��d�d�d�d�f�m�F��I����FǻN��E��e�e�d�e�g�l�F��H����V��_�E��y�_�u�u�g�m�G��H����V��_�D��d�e�e�d�f�m�[�ԜY���V��^�E��e�d�d�d�f�l�F��I����W�d��U���e�e�d�d�f�m�G��I����W��^�D��d�w�u�u�w��G��H����V��_�D��d�d�d�d�g�m�F���Y���D��^�E��e�e�e�d�g�l�F��H����V��L����u�e�e�e�g�l�G��H����W��_�E��d�e�d�y�]�}�W��I����W��^�D��e�d�d�d�f�m�F��H���F�^�E��d�d�e�e�g�l�F��H����W��_�W���u�u�w�e�g�l�F��I����V��_�D��e�d�d�e�u�}�W���[����W��_�E��d�d�e�d�f�l�F��H����FǻN��E��e�e�d�d�g�l�F��I����W��^�D��y�_�u�u�g�m�G��H����W��^�E��e�e�e�e�f�m�[�ԜY���V��^�D��e�e�d�e�g�m�G��H����V�d��U���e�e�d�d�f�m�F��I����V��^�D��e�w�u�u�w��G��H����V��_�D��e�e�e�d�f�m�F���Y���D��^�E��d�e�e�d�f�l�G��I����V��L����u�e�e�e�g�l�G��I����W��^�D��e�e�e�y�]�}�W��I����W��_�E��e�e�e�e�f�m�F��I���F�^�E��d�d�e�e�f�m�G��I����W��_�W���u�u�w�e�g�l�F��H����V��^�E��d�e�d�d�u�}�W���[����W��^�E��d�d�d�e�g�m�F��I����FǻN��E��e�e�d�e�g�l�F��H����W��^�D��y�_�u�u�g�m�G��H����W��_�E��e�e�e�d�f�l�[�ԜY���V��^�D��e�e�d�d�g�m�G��H����W�d��U���e�e�d�d�f�l�F��H����V��^�E��e�w�u�u�w��G��H����V��_�E��e�e�d�d�g�l�F���Y���D��^�E��d�d�d�d�g�m�G��H����W��L����u�e�e�e�g�m�G��H����W��^�D��d�e�e�y�]�}�W��I����W��_�D��e�e�e�e�f�l�G��H���F�^�E��e�d�d�d�g�l�F��I����V��^�W���u�u�w�e�g�l�G��I����W��^�E��d�e�e�d�u�}�W���[����W��^�E��d�d�e�e�g�l�F��I����FǻN��E��e�e�e�d�f�l�F��I����V��_�E��y�_�u�u�g�m�G��I����V��_�E��d�e�d�e�f�m�[�ԜY���V��^�E��e�d�e�d�g�m�F��H����W�d��U���e�e�d�e�g�l�F��H����V��^�D��d�w�u�u�w��G��I����V��_�E��e�e�e�d�g�m�F���Y���D��^�D��e�e�e�d�g�l�G��I����W��L����u�e�e�e�f�l�G��I����W��^�D��e�e�e�y�]�}�W��I����V��^�E��d�e�e�d�f�l�F��H���F�^�E��d�d�e�d�g�l�G��I����W��^�W���u�u�w�e�g�m�F��H����W��^�E��d�d�e�e�u�}�W���[����V��_�D��e�d�e�e�g�m�F��I����FǻN��E��e�d�d�d�f�l�F��I����V��_�E��y�_�u�u�g�m�G��H����W��_�E��d�e�e�e�f�l�[�ԜY���V��_�D��e�d�d�d�g�m�F��I����W�d��U���e�e�e�e�g�m�F��H����V��^�E��e�w�u�u�w��G��I����W��_�D��e�e�d�e�f�l�F���Y���D��^�E��d�d�d�d�g�l�G��H����W��L����u�e�e�e�g�l�G��H����W��^�E��e�e�e�y�]�}�W��I����V��^�E��d�e�e�d�g�l�G��H���F�^�E��d�e�d�d�f�m�F��I����W��_�W���u�u�w�e�g�m�G��I����W��^�E��d�d�e�d�u�}�W���[����V��^�D��d�d�d�e�g�l�G��H����FǻN��E��e�e�e�d�g�l�F��I����W��_�E��y�_�u�u�g�m�G��I����W��_�E��d�d�e�d�f�l�[�ԜY���V��^�E��e�e�e�e�g�m�F��H����W�d��U���d�d�d�d�f�m�F��H����V��_�E��d�w�u�u�w��F��H����V��^�D��e�e�d�e�f�m�G���Y���D��_�D��e�d�d�d�f�m�G��H����V��L����u�d�d�d�f�m�G��H����V��^�D��d�e�d�y�]�}�W��H����W��^�E��e�e�e�d�f�m�G��I���F�_�D��e�e�d�e�g�l�G��I����V��^�W���u�u�w�d�f�l�G��H����W��^�E��d�e�e�e�u�}�W���[����W��^�E��e�d�d�e�g�l�F��I����FǻN��D��d�e�d�d�g�m�F��H����W��^�D��y�_�u�u�f�l�F��H����V��^�E��d�d�e�d�g�l�[�ԜY���W��^�D��e�d�e�e�g�m�F��I����V�d��U���d�d�d�d�g�m�F��I����V��_�E��d�w�u�u�w��F��H����W��_�E��e�e�d�d�g�m�G���Y���D��_�E��d�e�d�e�f�l�G��H����W��L����u�d�d�d�g�m�F��H����W��^�D��d�e�d�y�]�}�W��H����V��^�E��e�e�e�d�f�l�G��I���F�_�D��e�e�e�d�f�l�F��I����W��_�W���u�u�w�d�f�m�F��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�d�d�e�g�l�G��I����FǻN��D��d�d�e�e�f�m�G��I����W��^�D��y�_�u�u�f�l�F��I����V��^�E��d�d�e�e�f�m�[�ԜY���W��_�D��e�d�e�e�g�m�F��H����W�d��U���d�d�e�e�g�l�G��I����V��^�E��d�w�u�u�w��F��I����W��_�D��e�e�d�d�f�m�F���Y���D��_�D��e�d�e�d�f�l�G��H����V��L����u�d�d�d�f�m�G��I����W��^�E��d�d�e�y�]�}�W��H����W��^�E��d�e�e�d�g�l�F��I���F�_�D��d�e�d�e�g�l�G��I����V��_�W���u�u�w�d�f�m�F��I����V��^�E��e�e�d�e�u�}�W���[����V��_�E��d�e�d�e�g�m�F��I����FǻN��D��d�e�e�d�g�l�F��I����V��_�D��y�_�u�u�f�l�F��H����W��^�E��d�d�e�e�g�m�[�ԜY���W��^�D��d�e�e�e�g�m�F��H����W�d��U���d�d�e�e�g�m�G��H����V��_�D��e�w�u�u�w��F��I����W��_�D��e�e�e�d�f�l�G���Y���D��_�E��e�e�e�e�f�m�G��I����W��L����u�d�d�d�g�m�F��I����V��^�E��d�d�e�y�]�}�W��H����V��_�D��d�e�e�d�g�l�F��I���F�_�D��d�d�e�d�g�l�G��I����V��_�W���u�u�w�d�f�l�F��I����V��^�E��d�d�d�e�u�}�W���[����W��^�D��e�d�e�e�g�l�F��I����FǻN��D��e�d�d�e�g�l�F��H����W��_�D��y�_�u�u�f�l�G��I����W��^�E��e�d�e�d�f�l�[�ԜY���W��_�D��e�e�d�e�g�m�G��H����V�d��U���d�d�d�d�f�m�F��I����V��^�D��e�w�u�u�w��F��H����W��^�E��e�e�d�e�f�m�F���Y���D��_�D��d�e�d�e�g�m�G��H����V��L����u�d�d�e�f�m�G��H����V��^�D��e�d�d�y�]�}�W��H����V��_�E��d�e�e�e�f�m�G��I���F�_�D��e�d�d�d�f�l�F��I����W��_�W���u�u�w�d�f�l�G��H����W��^�E��e�e�d�e�u�}�W���[����W��_�D��d�e�d�e�g�m�F��I����FǻN��D��e�d�d�d�f�l�G��H����V��^�D��y�_�u�u�f�l�G��H����V��^�E��e�e�d�e�g�m�[�ԜY���W��_�D��e�d�e�d�f�l�F��H����V�d��U���d�d�d�e�f�m�F��I����W��_�D��e�w�u�u�w��F��H����W��_�D��d�d�d�e�f�m�G���Y���D��_�D��d�d�e�e�f�l�F��H����V��L����u�d�d�e�f�m�G��H����V��_�E��e�e�d�y�]�}�W��H����V��_�E��d�d�d�d�g�l�F��I���F�_�D��d�e�d�d�g�l�F��H����V��_�W���u�u�w�d�f�l�F��I����W��_�D��d�d�e�e�u�}�W���[����W��_�E��e�d�e�d�f�m�F��I����FǻN��D��e�d�e�e�g�l�F��H����V��^�D��y�_�u�u�f�l�G��I����W��_�D��d�e�d�d�g�l�[�ԜY���W��_�E��e�d�d�d�f�l�F��I����W�d��U���d�d�d�d�g�m�F��H����W��^�E��d�w�u�u�w��F��H����V��^�D��d�d�e�e�g�m�G���Y���D��_�D��d�d�e�e�g�m�F��H����V��L����u�d�d�d�g�m�G��I����V��_�D��d�e�e�y�]�}�W��H����V��^�D��e�d�d�e�f�m�G��I���F�_�D��e�d�d�d�g�m�F��H����W��^�W���u�u�w�d�f�m�G��I����W��_�D��d�e�e�d�u�}�W���[����V��^�E��e�e�d�d�f�l�G��H����FǻN��D��d�e�d�d�g�m�F��I����W��^�E��y�_�u�u�f�l�F��I����W��_�D��e�d�e�d�g�l�[�ԜY���W��^�D��e�d�e�e�f�l�G��H����W�d��U���d�d�e�d�g�m�G��I����W��_�D��e�w�u�u�w��F��I����W��^�D��d�d�e�d�f�l�G���Y���D��_�E��d�e�e�d�g�m�F��I����V��L����u�d�d�d�f�m�F��H����W��_�E��e�e�d�y�]�}�W��H����V��^�D��e�d�d�e�g�m�G��I���F�_�D��e�e�d�e�g�l�G��H����W��^�W���u�u�w�d�f�m�G��H����V��_�E��d�d�e�e�u�}�W���[����V��^�D��d�e�d�d�g�l�G��I����FǻN��D��d�d�d�e�g�m�G��I����W��_�E��y�_�u�u�f�l�F��H����V��^�D��d�e�d�e�f�l�[�ԜY���W��^�E��d�e�e�d�f�l�F��I����V�d��U���d�d�d�e�f�m�G��I����W��^�E��d�w�u�u�w��F��H����V��_�E��d�e�d�e�g�l�F���Y���D��_�E��d�d�e�d�g�m�F��H����W��L����u�d�d�d�g�m�G��I����V��^�D��e�d�e�y�]�}�W��H����W��_�D��d�d�d�d�f�m�F��I���F�_�D��d�d�d�e�g�l�G��H����V��^�W���u�u�w�d�f�l�G��I����V��_�E��e�d�d�e�u�}�W���[����W��^�D��d�e�d�d�g�m�G��I����FǻN��D��d�d�d�d�g�m�F��I����V��^�D��y�_�u�u�f�l�F��I����V��^�D��d�e�d�d�g�l�[�ԜY���W��_�E��d�d�d�d�f�l�F��H����W�d��U���e�e�e�e�g�m�G��I����W��^�D��d�w�u�u�w��G��I����W��^�D��d�e�e�d�f�m�F���Y���D��^�E��d�e�d�d�g�l�F��I����W��L����u�e�e�e�g�m�G��H����V��^�E��d�d�e�y�]�}�W��I����V��_�D��e�d�d�d�g�l�G��H���F�^�E��d�d�e�d�f�m�G��H����W��_�W���u�u�w�e�g�m�G��I����W��_�E��e�e�e�d�u�}�W���[����V��^�D��e�e�e�d�g�m�G��H����FǻN��E��e�d�d�d�g�l�G��I����V��_�D��y�_�u�u�g�m�G��I����V��^�D��d�e�e�d�g�l�[�ԜY���V��_�E��d�e�d�e�f�l�F��I����V�d��U���e�e�d�e�g�m�G��H����W��^�D��e�w�u�u�w��G��H����V��_�D��d�e�e�e�f�m�F���Y���D��^�E��d�d�d�e�f�l�F��I����W��L����u�e�e�e�g�m�G��I����W��^�E��e�e�e�y�]�}�W��I����V��_�E��e�d�d�d�g�l�F��I���F�^�E��d�d�d�d�f�m�F��H����W��_�W���u�u�w�e�g�l�G��H����W��_�E��e�d�d�d�u�}�W���[����W��^�D��d�d�e�d�g�m�F��I����FǻN��E��e�d�d�d�f�m�G��I����V��_�D��y�_�u�u�g�m�G��I����W��^�D��d�e�d�e�g�l�[�ԜY���V��_�E��e�d�e�d�f�l�F��H����V�d��U���e�e�d�d�f�l�G��H����W��_�E��e�w�u�u�w��G��I����V��_�D��d�e�e�e�f�m�G���Y���D��^�E��e�d�d�d�f�l�F��I����W��L����u�e�e�d�g�l�F��H����V��^�D��e�e�d�y�]�}�W��I����V��^�E��d�d�d�d�f�m�F��H���F�^�E��d�e�d�d�f�m�G��H����W��_�W���u�u�w�e�g�m�F��I����V��_�E��e�d�e�e�u�}�W���[����V��^�E��e�d�e�d�g�l�G��H����FǻN��E��d�d�e�d�f�m�G��H����W��^�E��y�_�u�u�g�m�F��H����V��_�D��d�e�d�d�g�m�[�ԜY���V��_�E��d�e�d�d�f�l�F��I����V�d��U���e�e�e�d�f�l�G��H����W��_�E��d�w�u�u�w��G��I����W��^�D��d�e�d�d�f�m�F���Y���D��^�D��e�e�e�e�f�l�F��H����V��L����u�e�e�d�g�m�G��H����V��_�E��d�d�e�y�]�}�W��I����V��_�E��d�d�d�e�g�m�G��I���F�^�E��e�e�e�d�f�l�F��H����W��^�W���u�u�w�e�g�l�G��H����V��_�D��e�d�e�e�u�}�W���[����W��_�E��d�d�d�d�f�m�F��H����FǻN��E��d�e�e�d�g�l�F��I����V��_�D��y�_�u�u�g�m�F��I����V��_�D��e�e�d�e�f�m�[�ԜY���V��^�D��e�d�d�e�f�l�G��I����W�d��U���e�e�d�d�g�m�G��I����W��_�E��e�w�u�u�w��G��H����V��_�E��d�d�d�e�f�l�G���Y���D��^�E��d�d�e�e�f�m�F��H����W��L����u�e�e�d�f�m�G��H����V��_�E��d�d�e�y�]�}�W��I����V��^�E��e�d�d�d�g�m�G��I���F�^�E��e�e�d�e�g�l�G��H����V��^�W���u�u�w�e�g�l�G��I����V��_�D��e�d�d�e�u�}�W���[����W��_�D��e�d�e�d�f�m�F��H����FǻN��E��d�d�e�d�f�m�F��H����W��^�E��y�_�u�u�g�m�F��I����W��_�D��d�e�d�e�f�m�[�ԜY���V��_�D��d�e�e�d�f�l�F��H����V�d��U���e�e�d�e�f�l�F��I����W��_�D��e�w�u�u�w��G��H����W��_�D��e�e�e�e�f�l�G���Y���D��^�D��d�d�e�e�g�l�G��I����V��L����u�e�e�d�f�m�F��H����V��^�D��d�d�e�y�]�}�W��I����V��^�E��e�e�e�e�f�m�F��I���F�^�E��e�d�d�e�f�l�F��I����V��^�W���u�u�w�e�g�l�G��H����V��^�E��d�e�d�e�u�}�W���[����W��^�E��e�e�e�e�g�l�G��H����FǻN��E��d�d�e�e�f�m�G��I����W��^�D��y�_�u�u�g�m�F��H����V��^�E��d�e�e�e�g�m�[�ԜY���V��^�D��d�d�e�d�g�m�F��I����V�d��U���e�e�d�d�g�l�F��I����V��^�D��e�w�u�u�w��G��H����W��_�E��e�e�e�e�f�l�F���Y���D��^�E��e�e�e�d�g�l�G��I����W��L����u�e�e�d�g�m�G��I����W��^�E��d�d�e�y�]�}�W��I����W��^�E��d�e�e�d�g�l�F��H���F�^�E��e�e�d�e�g�m�F��I����W��^�W���u�u�w�e�g�l�G��H����W��^�E��d�d�d�e�u�}�W���[����W��^�D��e�e�d�e�f�m�G��H����FǻN��E��d�d�d�e�g�m�G��I����V��_�E��y�_�u�u�g�m�F��H����W��^�E��e�d�d�d�f�l�[�ԜY���V��_�E��d�d�d�d�g�m�G��H����V�d��U���e�e�e�e�f�m�F��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�d�d�d�g�m�G���Y���D��^�D��d�e�e�e�f�m�G��H����W��L����u�e�e�d�g�l�G��H����W��_�D��e�d�d�y�]�}�W��I����V��^�E��e�e�e�d�g�m�F��H���F�^�E��d�e�d�e�g�l�F��I����V��_�W���u�u�w�e�g�m�G��I����W��^�D��d�d�d�e�u�}�W���[����V��^�D��e�d�e�e�f�m�G��H����FǻN��E��e�d�d�e�g�m�F��I����V��^�E��y�_�u�u�g�m�G��I����W��_�E��d�e�e�d�g�l�[�ԜY���V��_�D��e�d�e�e�g�m�F��I����W�d��U���e�e�d�e�f�l�G��I����V��_�E��e�w�u�u�w��G��H����W��^�D��e�d�d�e�f�m�G���Y���D��^�E��d�d�e�e�g�m�G��H����V��L����u�e�e�e�g�l�F��H����W��^�E��d�d�d�y�]�}�W��I����V��^�D��e�e�d�e�g�l�F��H���F�^�E��d�d�e�d�f�l�F��H����W��^�W���u�u�w�e�g�m�F��I����V��^�E��e�e�d�d�u�}�W���[����V��_�D��e�e�e�e�g�m�G��H����FǻN��E��e�d�e�e�f�l�F��I����V��_�D��y�_�u�u�g�m�G��H����W��^�E��e�d�d�d�f�m�[�ԜY���V��^�E��e�d�d�d�g�l�G��I����W�d��U���e�e�e�e�g�l�F��H����W��^�D��d�w�u�u�w��G��I����V��^�E��e�e�d�d�f�l�G���Y���D��_�D��d�d�e�e�f�m�G��H����V��L����u�d�d�d�f�l�G��H����V��^�D��e�e�e�y�]�}�W��H����V��^�E��e�e�d�e�f�l�F��I���F�_�D��d�e�d�e�g�m�F��H����V��_�W���u�u�w�d�f�l�G��H����W��^�E��d�d�d�e�u�}�W���[����W��_�D��e�d�e�e�g�l�F��H����FǻN��D��d�d�d�d�f�m�F��I����W��_�D��y�_�u�u�f�l�F��I����V��_�E��d�e�e�e�g�m�[�ԜY���W��_�D��e�d�e�d�g�l�F��I����V�d��U���d�d�e�d�f�l�G��H����W��^�D��d�w�u�u�w��F��I����W��^�D��e�e�e�e�f�l�G���Y���D��_�E��e�e�d�e�g�l�G��I����V��L����u�d�d�e�f�l�F��I����V��^�E��e�d�e�y�]�}�W��H����V��^�E��e�e�d�d�g�l�G��H���F�_�D��e�e�d�e�g�m�G��H����V��_�W���u�u�w�d�f�l�G��I����V��^�E��e�d�e�e�u�}�W���[����W��_�D��d�d�d�e�g�m�G��H����FǻN��D��e�e�d�e�f�m�G��H����V��^�D��y�_�u�u�f�l�G��I����W��_�E��e�d�d�e�f�m�[�ԜY���W��_�E��d�d�d�e�g�l�G��H����W�d��U���d�d�e�e�f�l�G��I����W��_�D��e�w�u�u�w��F��I����W��^�E��e�e�d�e�f�l�G���Y���D��_�E��d�d�e�d�g�l�G��H����W��L����u�d�d�e�g�m�F��I����W��^�D��d�e�e�y�]�}�W��H����W��_�D��d�e�d�e�g�l�F��H���F�_�E��d�d�d�e�g�m�G��H����V��_�W���u�u�w�d�g�l�F��I����V��^�E��e�e�e�e�u�}�W���[����W��_�E��e�e�e�e�g�l�G��I����FǻN��D��d�d�e�e�f�m�G��I����V��_�E��y�_�u�u�f�l�F��H����V��^�E��e�d�d�d�f�l�[�ԜY���W��^�E��d�d�e�e�g�l�G��I����W�d��U���d�e�d�e�g�l�G��I����W��^�D��e�w�u�u�w��F��H����V��^�D��e�e�e�e�f�l�F���Y���D��^�D��d�e�e�e�f�l�G��H����W��L����u�d�d�d�f�m�F��I����W��_�D��d�d�e�y�]�}�W��H����W��_�E��d�e�e�d�g�l�G��I���F�_�E��e�d�e�e�g�m�G��I����W��_�W���u�u�w�d�g�m�F��H����W��^�D��d�d�d�e�u�}�W���[����V��_�E��e�e�e�e�f�m�G��I����FǻN��D��d�e�e�e�f�m�G��I����V��^�D��y�_�u�u�f�l�F��H����W��^�E��d�e�d�e�f�l�[�ԜY���W��^�D��e�d�e�e�g�m�G��I����V�d��U���d�e�d�d�f�l�G��I����V��_�E��d�w�u�u�w��F��H����W��^�E��e�d�d�d�g�m�G���Y���D��^�D��e�d�e�e�f�m�G��I����W��L����u�d�d�e�f�m�G��H����V��_�D��d�d�e�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��I���F�_�E��e�e�e�e�g�l�G��I����W��^�W���u�u�w�d�g�l�G��I����W��^�E��e�d�e�e�u�}�W���[����W��^�E��d�d�e�e�g�l�G��H����FǻN��D��e�e�d�d�g�l�F��H����V��_�D��y�_�u�u�f�l�G��H����W��_�E��d�e�d�e�g�l�[�ԜY���W��^�E��d�e�e�d�g�m�F��I����W�d��U���d�e�d�d�g�m�G��I����V��_�E��d�w�u�u�w��F��H����V��^�E��e�e�d�d�g�l�G���Y���D��^�E��d�e�e�d�f�m�G��I����W��L����u�d�d�e�g�m�G��I����W��^�E��e�d�d�y�]�}�W��H����V��_�D��e�e�e�e�g�m�G��H���F�_�E��d�d�d�d�f�m�F��H����V��^�W���u�u�w�d�g�l�F��I����V��_�D��e�e�e�e�u�}�W���[����W��^�E��d�e�e�d�f�m�G��I����FǻN��D��e�e�d�e�f�m�G��H����V��^�D��y�_�u�u�f�l�G��H����W��_�D��e�d�e�e�f�l�[�ԜY���W��^�D��e�e�e�d�f�l�G��I����W�d��U���d�e�d�e�g�l�G��I����W��_�E��d�w�u�u�w��F��H����W��^�D��d�d�e�d�g�l�F���Y���D��^�D��e�e�e�e�g�m�F��H����W��L����u�d�d�e�f�l�G��I����V��^�E��d�e�e�y�]�}�W��H����V��_�D��d�d�d�d�g�m�G��H���F�_�E��d�e�e�d�g�l�G��H����V��_�W���u�u�w�d�g�l�F��I����W��_�E��e�e�e�e�u�}�W���[����V��_�D��e�d�d�d�g�l�G��H����FǻN��D��d�e�d�d�f�l�G��H����W��^�D��y�_�u�u�f�l�F��I����V��^�D��e�d�e�e�g�l�[�ԜY���W��^�E��e�e�e�e�f�l�G��I����V�d��U���d�e�e�e�g�l�F��H����V��_�D��e�w�u�u�w��F��I����V��_�D��d�d�d�e�f�l�G���Y���D��^�D��e�d�e�e�g�l�F��I����W��L����u�d�d�d�f�l�F��H����V��_�E��e�e�d�y�]�}�W��H����W��^�D��d�d�e�e�f�m�G��I���F�_�E��d�d�d�e�g�m�F��I����V��_�W���u�u�w�d�g�l�G��I����W��_�D��e�d�d�d�u�}�W���[����W��_�E��e�e�e�d�f�m�G��I����FǻN��D��d�d�d�e�f�l�F��H����W��_�E��y�_�u�u�f�l�G��I����V��_�D��d�e�e�d�f�m�[�ԜY���W��^�E��e�e�e�e�f�m�F��I����V�d��U���d�d�e�e�g�m�F��I����V��^�E��e�w�u�u�w��F��I����W��_�D��d�e�d�e�g�m�F���Y���D��_�D��d�e�e�e�f�m�F��H����V��L����u�d�d�e�g�l�G��H����V��^�D��d�e�e�y�]�}�W��H����W��^�D��e�d�e�e�g�l�G��H���F�_�D��e�d�d�d�f�l�G��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��d�e�e�d�u�}�W���[����V��_�E��d�e�e�e�f�m�F��H����FǻN��D��d�d�e�e�g�m�G��I����V��_�E��y�_�u�u�f�l�F��I����W��_�D��e�d�d�e�g�l�[�ԜY���W��^�D��e�d�d�d�f�l�G��H����W�d��U���d�d�d�d�g�m�G��I����W��^�E��e�w�u�u�w��F��H����V��^�D��e�d�e�e�f�m�F���Y���D��^�E��e�e�e�e�g�m�G��I����W��L����u�e�e�e�g�m�G��I����V��^�D��d�e�e�y�]�}�W��I����W��_�D��d�d�d�d�g�m�G��I���F�^�E��d�d�e�e�g�l�F��H����W��^�W���u�u�w�e�g�l�F��H����W��_�E��e�e�d�d�u�}�W���[����W��^�E��d�e�d�e�g�m�G��H����FǻN��E��e�d�d�d�f�m�G��H����W��^�E��y�_�u�u�g�m�F��I����W��_�D��e�e�d�e�f�l�[�ԜY���V��_�D��e�e�d�e�f�l�G��I����V�d��U���e�e�d�e�f�m�F��I����W��_�D��e�w�u�u�w��G��H����V��_�D��e�e�e�d�f�m�F���Y���D��^�D��e�e�e�d�f�l�G��I����V��L����u�e�e�e�g�l�G��I����W��_�D��e�d�e�y�]�}�W��I����V��_�E��d�d�e�d�g�l�F��I���F�^�D��d�d�d�d�f�m�F��I����V��^�W���u�u�w�e�f�l�F��I����V��_�D��d�d�d�d�u�}�W���[����W��^�E��d�d�d�e�f�m�G��I����FǻN��E��d�e�d�d�g�m�F��I����V��^�D��y�_�u�u�g�m�F��I����V��_�D��d�e�e�d�f�m�[�ԜY���V��_�D��e�d�e�e�f�m�G��I����W�d��U���e�d�d�d�g�m�G��H����V��_�D��d�w�u�u�w��G��H����W��_�E��e�d�d�d�g�l�G���Y���D��^�E��d�e�e�e�g�l�G��H����W��L����u�e�d�e�f�l�G��I����V��_�E��e�e�d�y�]�}�W��H����V��^�E��d�d�e�e�f�m�F��I���F�^�E��d�d�d�d�f�m�G��I����W��_�W���u�u�w�e�g�l�F��I����V��_�D��e�e�d�d�u�}�W���[����V��_�E��e�d�d�e�f�m�F��H����FǻN��E��d�d�e�d�g�m�F��H����V��_�D��y�_�u�u�g�l�F��H����W��^�D��e�e�d�d�f�m�[�ԜY���W��_�E��d�e�e�e�f�m�G��H����V�d��U���e�d�e�e�f�l�G��H����V��^�D��d�w�u�u�w��G��I����W��^�D��e�d�e�e�g�l�G���Y���D��_�D��e�d�d�d�f�m�G��H����W��L����u�e�d�e�g�l�G��H����W��^�D��e�d�d�y�]�}�W��H����V��_�D��d�d�e�d�f�l�G��H���F�^�D��d�e�d�d�g�m�G��I����W��_�W���u�u�w�e�f�m�G��H����W��_�E��d�d�d�e�u�}�W���[����W��^�D��e�d�e�e�f�m�G��H����FǻN��E��d�d�e�e�f�l�G��H����V��_�D��y�_�u�u�g�m�G��I����V��^�D��e�e�d�e�g�m�[�ԜY���V��^�D��d�d�e�d�f�m�G��H����W�d��U���d�e�e�d�g�m�F��H����V��^�D��e�w�u�u�w��F��H����V��^�E��e�d�e�d�f�m�F���Y���D��^�D��d�d�d�d�f�l�G��I����V��L����u�e�e�d�g�l�F��I����W��_�D��d�e�e�y�]�}�W��I����V��^�E��d�d�e�e�f�l�G��H���F�^�E��e�e�d�d�f�m�F��I����V��_�W���u�u�w�d�g�l�F��I����V��_�D��e�d�d�d�u�}�W���[����W��_�D��d�d�e�e�f�l�F��H����FǻN��E��e�e�e�e�f�l�G��I����W��^�E��y�_�u�u�g�m�G��H����V��^�D��e�d�d�d�f�m�[�ԜY���V��^�D��d�d�d�d�f�m�F��H����W�d��U���d�d�d�d�f�m�F��H����V��^�E��d�w�u�u�w��F��H����W��_�D��e�d�e�e�f�l�F���Y���D��_�E��e�d�d�e�g�m�G��H����V��L����u�e�e�d�f�l�G��H����W��_�E��e�d�d�y�]�}�W��I����V��_�D��d�d�e�d�f�l�G��H���F�^�D��d�e�d�d�g�m�G��I����W��^�W���u�u�w�d�f�l�F��H����V��_�E��d�d�d�d�u�}�W���[����V��^�D��e�e�e�e�g�m�G��H����FǻN��E��e�e�d�d�f�m�F��H����W��_�D��y�_�u�u�g�l�G��I����W��_�D��e�e�d�d�f�l�[�ԜY���W��^�D��d�e�e�e�f�l�G��H����W�d��U���d�e�d�e�g�l�F��I����W��^�E��d�w�u�u�w��F��H����W��_�D��e�e�e�e�f�l�G���Y���D��^�E��e�e�e�e�f�m�G��H����V��L����u�e�d�d�f�m�G��I����V��^�D��e�d�e�y�]�}�W��H����V��^�D��d�d�d�e�g�m�F��I���F�^�E��e�d�d�e�g�l�G��H����V��^�W���u�u�w�d�g�l�F��I����W��_�D��e�d�e�e�u�}�W���[����W��_�D��e�d�d�e�f�l�G��I����FǻN��E��d�d�d�d�f�m�G��I����V��_�E��y�_�u�u�g�l�G��I����W��^�D��d�d�d�e�g�l�[�ԜY���W��_�E��e�e�e�e�f�l�F��H����V�d��U���d�d�e�d�g�l�F��I����W��_�D��e�w�u�u�w��F��H����V��_�D��d�e�e�d�g�m�G���Y���D��_�E��e�e�d�e�f�m�F��I����V��L����u�e�d�e�g�l�F��H����W��^�E��d�e�e�y�]�}�W��H����W��_�D��e�d�e�d�g�m�G��I���F�^�D��d�e�e�e�f�m�F��I����V��_�W���u�u�w�d�f�m�G��I����W��_�E��e�d�d�e�u�}�W���[����V��^�E��e�d�d�d�g�l�F��I����FǻN��E��d�e�d�d�f�l�F��H����V��^�D��y�_�u�u�g�l�F��H����V��_�D��e�e�e�d�g�l�[�ԜY���W��_�E��d�e�d�e�f�m�G��H����W�d��U���d�d�e�d�f�l�G��I����V��^�D��d�w�u�u�w��F��H����V��^�E��d�d�e�d�f�l�G���Y���D��_�E��d�e�e�d�g�l�F��H����V��L����u�e�d�d�g�m�F��I����V��^�E��e�d�d�y�]�}�W��H����W��_�D��e�d�d�e�f�l�F��I���F�^�D��e�d�e�d�g�m�G��H����V��^�W���u�u�w�d�f�l�G��I����V��_�E��e�d�d�e�u�}�W���[����W��_�E��d�d�d�d�g�m�F��I����FǻN��E��d�d�e�d�f�m�F��I����W��_�D��y�_�u�u�g�l�F��I����V��_�D��e�e�e�e�f�l�[�ԜY���W��_�E��d�d�d�d�f�l�G��H����V�d��U���d�d�d�d�f�m�G��I����W��_�D��d�w�u�u�w��F��H����V��^�D��d�d�e�d�g�m�F���Y���D��_�D��d�e�d�e�g�l�F��I����V��L����u�e�d�d�f�l�F��I����W��_�D��d�e�d�y�]�}�W��H����W��^�D��e�e�e�e�g�m�G��H���F�^�D��d�d�e�d�g�l�G��I����V��_�W���u�u�w�d�f�l�F��I����V��^�E��e�d�d�e�u�}�W���[����W��^�E��e�d�d�e�g�m�F��I����FǻN��E��d�d�e�d�g�m�G��H����W��_�E��y�_�u�u�g�l�F��I����V��_�E��d�d�d�d�g�l�[�ԜY���W��_�D��e�d�d�d�g�m�G��H����V�d��U���d�d�d�e�g�m�G��I����V��^�D��e�w�u�u�w��F��H����V��^�E��e�d�d�d�g�m�F���Y���D��_�E��e�d�e�d�g�m�G��I����W��L����u�e�d�d�g�m�F��I����V��_�E��e�e�e�y�]�}�W��H����W��^�E��d�e�e�d�f�l�F��H���F�^�D��e�d�e�e�g�l�F��H����W��^�W���u�u�w�d�f�m�F��H����V��^�E��e�e�e�e�u�}�W���[����V��^�D��d�e�d�e�g�l�G��H����FǻN��E��d�d�d�e�f�m�F��I����V��_�E��y�_�u�u�g�l�F��H����W��^�E��d�d�d�e�f�l�[�ԜY���W��^�E��e�d�d�e�g�l�F��I����V�d��U���d�d�e�e�f�m�F��H����W��^�E��d�w�u�u�w��F��H����V��_�D��e�d�e�d�g�m�F���Y���D��_�D��e�d�d�e�f�m�G��H����W��L����u�e�d�e�g�l�F��H����W��_�D��d�e�e�y�]�}�W��H����V��^�E��e�e�d�d�f�m�G��I���F�^�D��e�e�e�d�f�l�F��H����W��_�W���u�u�w�d�f�m�F��H����V��^�D��e�d�d�d�u�}�W���[����V��^�E��e�d�d�d�g�m�F��H����FǻN��E��e�e�e�e�g�l�G��H����V��_�D��y�_�u�u�g�l�F��H����V��^�E��e�e�e�d�f�l�[�ԜY���W��_�D��d�d�e�e�g�m�G��H����W�d��U���d�e�d�d�g�m�G��H����V��^�E��e�w�u�u�w��F��H����W��^�E��d�e�e�d�g�m�G���Y���D��^�D��e�e�d�d�g�l�F��H����W��L����u�e�d�d�f�m�G��I����V��^�D��e�d�e�y�]�}�W��H����W��^�E��e�e�e�e�g�m�F��I���F�^�E��d�d�d�e�f�m�G��I����V��_�W���u�u�w�d�g�l�G��H����V��^�D��d�e�e�d�u�}�W���[����W��_�E��e�e�e�d�f�l�G��I����FǻN��E��e�d�e�d�g�l�G��H����V��_�E��y�_�u�u�g�l�G��H����V��_�E��d�d�e�e�g�l�[�ԜY���W��^�E��e�d�d�d�g�m�F��H����W�d��U���d�d�d�d�g�l�F��I����V��^�E��d�w�u�u�w��F��H����W��^�E��d�d�d�e�g�m�F���Y���D��_�E��e�d�d�d�g�m�F��I����V��L����u�e�e�d�f�l�G��H����W��^�E��d�d�d�y�]�}�W��I����V��_�D��d�e�d�e�f�l�F��H���F�^�D��d�d�d�e�f�l�F��H����W��^�W���u�u�w�d�f�l�F��I����W��^�E��d�e�e�d�u�}�W���[����W��_�D��d�e�d�d�g�l�G��I����FǻN��E��e�d�d�d�g�m�F��I����W��_�E��y�_�u�u�g�m�G��I����W��_�E��d�e�e�e�f�m�[�ԜY���V��_�D��e�d�d�d�g�l�F��I����W�d��U���d�e�d�d�f�m�G��I����W��_�E��d�w�u�u�w��F��H����W��_�D��d�e�e�d�g�m�G���Y���D��^�D��d�e�d�e�g�l�F��I����V��L����u�e�e�d�g�l�F��I����W��^�E��d�d�d�y�]�}�W��I����W��_�D��e�e�d�d�g�m�F��I���F�^�E��d�d�e�e�g�l�F��H����W��^�W���u�u�w�d�g�m�F��I����W��^�E��e�e�d�e�u�}�W���[����V��_�E��e�d�e�d�g�l�G��H����FǻN��E��e�e�e�e�f�m�F��H����W��^�E��y�_�u�u�g�l�F��I����W��_�E��d�d�e�d�f�m�[�ԜY���W��^�E��d�e�d�e�g�l�F��H����W�d��U���e�d�e�e�f�l�F��H����W��_�D��e�w�u�u�w��G��I����W��^�E��d�d�e�e�g�l�G���Y���D��_�D��e�d�d�d�f�m�F��I����V��L����u�e�d�e�g�l�G��H����W��_�E��d�d�d�y�]�}�W��H����W��_�E��e�e�d�e�g�m�F��H���F�^�D��e�e�d�e�g�l�G��H����V��_�W���u�u�w�e�f�m�G��H����W��^�E��d�d�e�e�u�}�W���[����W��^�D��e�e�d�d�g�l�F��H����FǻN��E��d�e�d�e�f�l�G��H����W��_�D��y�_�u�u�g�l�F��I����V��_�E��d�d�e�e�f�m�[�ԜY���W��^�D��d�d�e�e�g�l�F��H����V�d��U���e�e�d�d�g�m�F��I����W��_�D��e�w�u�u�w��G��H����W��_�D��d�e�d�d�f�m�G���Y���D��^�E��e�e�d�e�g�l�F��H����W��L����u�e�d�e�f�l�G��I����V��^�E��e�e�e�y�]�}�W��H����W��^�E��d�e�d�d�f�l�F��H���F�^�D��d�e�d�e�f�m�F��H����V��^�W���u�u�w�e�f�l�F��I����W��^�E��e�d�e�e�u�}�W���[����V��_�E��d�d�d�d�g�m�F��H����FǻN��E��d�d�e�e�g�m�F��I����V��^�E��y�_�u�u�g�m�F��H����V��^�E��e�d�d�e�g�m�[�ԜY���V��_�E��d�e�e�d�g�l�G��H����V�d��U���e�d�d�d�f�m�F��I����W��^�E��d�w�u�u�w��G��I����W��_�E��d�e�d�e�g�m�G���Y���D��_�D��e�d�d�d�f�m�F��I����V��L����u�e�e�e�g�l�G��I����W��^�D��e�d�e�y�]�}�W��I����V��^�E��e�e�d�e�g�m�F��I���F�^�E��d�d�e�e�f�l�G��I����W��^�W���u�u�w�e�g�l�G��I����V��^�D��e�e�d�e�u�}�W���[����V��_�E��e�e�e�d�f�l�F��H����FǻN��E��d�e�e�d�g�l�F��I����V��_�E��y�_�u�u�g�m�G��H����V��^�E��d�d�e�d�g�l�[�ԜY���V��_�E��d�d�e�d�g�m�F��H����W�d��U���e�e�d�d�g�l�F��H����V��_�D��d�w�u�u�w��G��I����V��^�E��d�d�d�d�f�m�F���Y���D��^�D��e�d�d�e�g�m�F��H����W��L����u�e�e�e�g�m�G��I����V��_�D��d�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�_�D��e�d�e�e�g�l�F��I����V��^�W���u�u�w�d�f�l�F��I����V��^�E��d�e�d�e�u�}�W���[����W��_�D��d�e�e�d�g�m�F��H����FǻN��D��d�d�e�d�g�l�F��H����V��^�E��y�_�u�u�f�l�F��I����V��^�E��d�e�e�d�f�l�[�ԜY���W��^�D��d�e�d�e�g�m�G��H����V�d��U���d�d�d�d�f�m�G��I����V��^�D��d�w�u�u�w��F��H����W��_�E��d�e�e�e�f�l�F���Y���D��_�E��e�e�d�e�f�l�F��I����W��L����u�d�d�e�g�l�G��H����V��_�D��d�e�d�y�]�}�W��H����W��^�D��d�e�d�d�g�m�G��I���F�_�D��e�d�d�e�f�l�F��H����V��^�W���u�u�w�d�f�m�G��I����V��^�D��d�d�d�e�u�}�W���[����V��^�E��e�d�d�e�f�l�F��I����FǻN��D��e�e�e�e�f�m�F��H����W��^�D��y�_�u�u�f�l�F��H����W��_�E��e�d�d�e�g�m�[�ԜY���W��_�D��d�d�d�e�g�l�G��H����V�d��U���d�e�d�e�g�m�F��H����W��_�E��e�w�u�u�w��F��H����W��^�D��e�e�d�d�g�m�F���Y���D��^�E��d�e�e�d�g�m�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��d�d�e�y�]�}�W��H����V��_�E��e�e�d�e�f�l�F��H���F�_�E��e�d�e�d�f�m�G��H����W��_�W���u�u�w�d�g�m�G��H����W��^�E��d�e�e�d�u�}�W���[����V��^�E��e�d�d�e�g�m�F��H����FǻN��D��d�e�e�d�g�m�G��I����W��^�E��y�_�u�u�f�l�F��H����W��_�E��d�e�d�d�f�l�[�ԜY���W��^�D��e�d�d�e�g�m�F��H����W�d��U���d�e�d�d�f�m�F��H����V��^�D��e�w�u�u�w��F��H����V��^�D��e�d�d�d�f�l�F���Y���D��^�D��d�d�e�e�g�m�G��H����V��L����u�d�d�e�f�l�G��I����V��_�D��d�e�d�y�]�}�W��H����W��^�D��e�e�e�e�f�m�G��I���F�_�E��e�d�d�d�g�m�F��I����V��^�W���u�u�w�d�g�l�G��H����V��^�E��e�d�e�e�u�}�W���[����W��_�D��e�e�d�e�g�l�G��I����FǻN��D��e�e�d�d�f�l�F��H����V��^�D��y�_�u�u�f�l�G��H����V��^�E��d�e�d�d�g�l�[�ԜY���W��^�E��e�d�e�e�g�m�G��H����W�d��U���d�e�d�d�f�m�F��I����V��^�E��d�w�u�u�w��F��H����W��_�D��e�e�e�d�f�l�G���Y���D��^�E��e�d�e�e�g�m�G��I����W��L����u�d�d�e�g�m�G��I����W��_�D��d�e�d�y�]�}�W��H����V��^�E��d�d�d�d�f�m�F��H���F�_�E��d�d�e�d�g�l�F��H����W��_�W���u�u�w�d�g�l�F��I����V��_�D��e�d�e�d�u�}�W���[����W��^�D��e�e�e�d�f�m�F��I����FǻN��D��e�e�d�d�f�l�G��I����W��^�E��y�_�u�u�f�l�G��H����W��^�D��e�d�e�d�f�l�[�ԜY���W��_�E��e�d�d�d�f�l�G��H����W�d��U���d�e�d�e�f�m�F��H����W��_�E��d�w�u�u�w��F��H����V��^�D��d�d�e�d�g�l�G���Y���D��^�D��d�d�d�e�f�l�F��I����V��L����u�d�d�e�f�m�G��H����V��^�D��d�d�e�y�]�}�W��H����V��_�D��e�d�d�d�g�l�G��I���F�_�E��d�e�d�d�g�m�F��H����V��^�W���u�u�w�d�g�l�F��H����V��_�E��e�d�d�d�u�}�W���[����V��_�D��e�e�d�d�g�m�F��I����FǻN��D��d�e�d�d�g�l�F��H����V��^�E��y�_�u�u�f�l�F��I����V��_�D��e�d�e�d�g�l�[�ԜY���W��^�D��e�e�e�d�f�l�G��I����V�d��U���d�e�e�d�f�l�G��H����W��^�E��e�w�u�u�w��F��I����V��^�D��d�e�d�e�g�m�G���Y���D��^�D��d�d�d�e�g�m�F��I����V��L����u�d�d�d�f�m�F��I����W��^�D��d�e�e�y�]�}�W��H����W��^�E��d�d�d�e�g�m�G��I���F�_�E��e�e�e�d�g�m�F��H����V��^�W���u�u�w�d�g�l�G��H����V��_�D��d�e�e�d�u�}�W���[����W��^�E��d�e�e�d�f�l�G��I����FǻN��D��d�e�d�d�f�m�F��I����W��_�D��y�_�u�u�f�l�F��I����V��_�D��d�e�e�e�g�l�[�ԜY���W��_�D��d�e�e�d�f�m�F��H����W�d��U���d�e�d�d�f�m�F��I����V��_�D��e�w�u�u�w��F��H����W��^�D��d�d�e�d�f�m�G���Y���D��_�E��e�d�e�e�g�l�F��I����W��L����u�d�d�e�g�m�F��I����W��_�D��e�e�d�y�]�}�W��H����W��_�E��d�d�e�d�g�l�G��I���F�_�D��e�d�d�d�g�l�F��I����V��^�W���u�u�w�d�f�m�G��H����V��_�D��d�e�e�d�u�}�W���[����V��^�D��d�e�d�d�f�m�G��H����FǻN��D��e�e�e�d�f�l�G��I����V��_�D��y�_�u�u�f�l�G��H����V��_�D��d�e�e�d�f�m�[�ԜY���W��^�D��d�d�e�d�f�m�G��H����W�d��U���d�d�d�e�g�m�F��I����V��_�D��d�w�u�u�w��F��H����W��^�D��d�d�d�d�g�m�G���Y���D��_�D��e�e�d�e�g�m�F��H����V��L����u�d�d�e�f�l�F��I����V��_�D��d�d�d�y�]�}�W��H����W��^�E��e�d�e�e�f�m�F��I���F�_�D��d�e�d�e�g�l�G��I����V��_�W���u�u�w�d�f�m�F��H����W��_�D��d�e�e�e�u�}�W���[����V��_�D��d�d�d�d�f�l�F��I����FǻN��D��d�d�e�e�f�m�F��H����W��_�E��y�_�u�u�f�l�F��H����V��_�D��e�d�d�d�g�m�[�ԜY���W��^�D��d�e�d�e�f�m�F��I����V�d��U���d�d�d�e�f�l�G��H����V��^�D��e�w�u�u�w��F��H����W��^�D��d�d�e�e�g�m�G���Y���D��_�D��d�e�e�e�f�m�F��I����W��L����u�d�d�d�f�l�G��H����V��_�E��e�e�e�y�]�}�W��H����V��_�E��e�d�e�d�g�l�F��I���F�^�E��e�e�e�e�g�m�G��I����V��_�W���u�u�w�e�g�m�G��H����W��_�D��e�e�e�e�u�}�W���[����V��^�D��d�e�d�d�f�m�F��I����FǻN��E��e�e�d�d�f�l�F��I����V��^�E��y�_�u�u�g�m�G��I����W��_�D��d�e�e�e�f�m�[�ԜY���V��_�D��e�d�d�d�f�m�F��H����V�d��U���e�e�e�d�f�m�F��I����V��^�E��d�w�u�u�w��G��I����V��_�D��d�d�d�d�f�m�G���Y���D��^�E��d�e�d�d�g�m�F��H����V��L����u�e�e�e�g�l�F��H����W��_�D��e�e�d�y�]�}�W��I����V��_�E��d�d�e�d�f�l�G��H���F�^�E��d�d�d�d�g�l�G��H����V��_�W���u�u�w�e�g�l�G��H����V��_�E��d�e�d�e�u�}�W���[����W��_�D��d�d�e�d�g�m�F��H����FǻN��E��e�d�e�e�f�l�F��H����V��^�D��y�_�u�u�g�m�G��H����V��^�D��e�d�d�e�f�l�[�ԜY���V��^�E��d�d�e�e�f�l�G��I����W�d��U���e�e�e�e�g�m�G��H����W��^�E��d�w�u�u�w��G��I����W��^�E��d�e�d�e�g�m�F���Y���D��^�E��d�e�d�d�g�l�F��H����V��L����u�e�e�d�g�l�G��H����W��^�D��e�e�d�y�]�}�W��I����V��^�D��e�d�d�d�g�l�F��H���F�^�E��e�e�e�d�g�l�G��H����W��_�W���u�u�w�e�g�m�G��I����V��_�E��e�d�d�e�u�}�W���[����V��^�E��e�d�e�d�g�m�F��I����FǻN��E��d�d�d�e�g�l�G��H����W��_�E��y�_�u�u�g�m�F��H����V��^�D��d�e�e�e�g�l�[�ԜY���V��^�E��e�e�e�d�f�l�F��I����W�d��U���e�e�d�e�f�l�G��H����W��_�E��e�w�u�u�w��G��H����W��^�D��d�d�e�e�g�m�G���Y���D��^�E��e�e�d�e�f�l�F��I����V��L����u�e�e�d�g�m�G��I����W��_�D��e�d�d�y�]�}�W��I����V��^�D��e�d�d�e�f�m�G��I���F�^�E��d�d�d�e�f�l�F��H����V��_�W���u�u�w�e�g�l�F��H����V��_�D��d�e�e�e�u�}�W���[����W��_�E��e�e�e�d�f�l�G��I����FǻN��E��d�e�d�d�f�m�G��I����W��^�E��y�_�u�u�g�m�F��I����V��_�D��e�d�d�d�f�m�[�ԜY���V��_�E��d�d�d�d�f�l�F��H����W�d��U���e�e�d�e�g�l�F��I����W��^�D��d�w�u�u�w��G��H����W��_�D��d�d�e�e�f�m�F���Y���D��^�D��d�e�d�d�g�m�F��I����W��L����u�e�e�d�f�m�F��H����V��_�E��e�e�e�y�]�}�W��I����V��_�E��d�d�d�d�g�l�G��I���F�^�E��e�d�d�d�f�m�F��H����W��_�W���u�u�w�e�g�l�G��H����V��_�D��d�e�e�e�u�}�W���[����W��_�D��e�d�d�e�g�m�G��H����FǻN��E��d�d�e�d�g�l�G��H����V��^�E��y�_�u�u�g�m�F��I����V��^�E��e�d�e�d�f�m�[�ԜY���V��_�D��d�d�d�e�g�m�G��I����W�d��U���e�e�d�e�f�m�F��I����V��^�E��e�w�u�u�w��G��H����W��^�D��e�e�d�d�g�m�F���Y���D��^�D��d�e�d�d�g�m�G��H����V��L����u�e�e�d�f�m�G��H����V��^�D��e�e�e�y�]�}�W��I����W��_�D��d�e�e�e�f�l�G��I���F�^�E��d�d�e�d�f�l�F��I����V��^�W���u�u�w�e�g�l�F��I����V��^�E��d�e�d�e�u�}�W���[����W��_�D��e�e�e�e�g�m�F��H����FǻN��E��d�e�e�e�g�m�G��I����V��^�D��y�_�u�u�g�m�F��I����W��^�E��d�d�e�d�f�m�[�ԜY���V��^�D��e�d�e�d�g�m�F��I����W�d��U���e�e�d�e�g�l�F��I����V��^�D��d�w�u�u�w��G��H����V��_�E��e�e�d�d�g�l�F���Y���D��^�E��e�d�d�d�g�m�G��H����V��L����u�e�e�d�g�m�G��H����V��^�D��d�e�e�y�]�}�W��I����W��^�D��e�e�e�d�f�l�G��I���F�^�E��d�e�d�d�g�m�F��I����V��^�W���u�u�w�e�g�m�F��H����W��^�D��e�e�d�d�u�}�W���[����V��^�D��d�e�e�e�f�m�F��I����FǻN��E��d�d�d�e�g�m�F��I����V��_�D��y�_�u�u�g�m�F��I����V��^�E��e�d�e�e�g�m�[�ԜY���V��_�E��e�d�e�e�g�m�G��H����W�d��U���e�e�e�d�f�m�F��I����V��_�D��d�w�u�u�w��G��I����W��_�D��e�d�e�d�g�l�G���Y���D��^�E��e�e�e�d�g�m�G��H����V��L����u�e�e�d�g�l�F��H����V��_�E��e�d�d�y�]�}�W��I����W��_�E��d�e�e�e�g�l�F��H���F�^�E��e�d�e�e�f�m�G��I����V��^�W���u�u�w�e�g�l�F��H����W��^�D��d�e�d�e�u�}�W���[����W��^�D��d�d�e�e�f�l�F��I����FǻN��E��e�d�e�e�g�l�G��I����W��^�D��y�_�u�u�g�m�G��H����V��^�E��e�d�e�d�f�l�[�ԜY���V��_�E��d�e�e�d�g�m�G��H����V�d��U���e�e�d�e�g�l�G��H����V��_�D��d�w�u�u�w��G��H����W��_�E��e�d�d�d�g�m�G���Y���D��^�E��d�d�d�e�g�l�G��H����W��L����u�e�e�e�g�m�G��I����W��_�D��e�e�e�y�]�}�W��I����W��_�D��d�e�e�e�f�m�F��I���F�^�E��e�d�e�e�f�m�G��I����W��^�W���u�u�w�e�g�l�G��I����W��^�D��d�e�d�d�u�}�W���[����V��^�E��e�d�e�e�f�l�F��H����FǻN��E��e�d�e�e�g�m�F��H����W��^�E��y�_�u�u�g�m�G��H����W��_�E��e�d�d�e�f�l�[�ԜY���V��_�E��e�d�e�d�g�m�G��H����W�d��U���e�e�e�e�g�m�G��H����V��_�E��e�w�u�u�w��G��I����V��_�D��e�d�d�d�f�l�G���Y���D��^�E��d�d�d�d�g�m�G��H����W��L����u�e�e�e�g�m�G��H����V��_�D��d�d�d�y�]�}�W��I����W��^�E��e�e�e�e�f�m�G��I���F�^�E��e�d�d�e�g�l�G��I����W��_�W���u�u�w�e�g�m�G��I����V��^�D��e�e�d�e�u�}�W���[����W��^�E��d�d�e�e�f�l�G��I����FǻN��D��d�d�e�e�f�m�F��H����W��_�D��y�_�u�u�f�l�F��H����V��_�E��e�d�e�e�f�l�[�ԜY���W��_�E��d�d�e�e�g�m�G��H����W�d��U���d�d�d�e�f�m�F��I����V��^�D��d�w�u�u�w��F��H����W��^�D��e�d�d�d�g�m�F���Y���D��_�E��e�d�d�e�f�m�G��H����W��L����u�d�d�d�g�m�G��I����V��_�E��e�e�e�y�]�}�W��H����W��_�E��e�e�e�e�g�m�F��I���F�_�D��e�e�e�d�f�m�F��I����W��_�W���u�u�w�d�f�l�G��I����V��^�D��d�d�e�d�u�}�W���[����W��^�E��e�e�d�e�f�m�G��H����FǻN��D��d�d�d�e�f�m�F��I����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�d�e�d�g�l�[�ԜY���W��_�E��e�e�e�d�g�m�G��H����W�d��U���d�d�e�e�f�l�F��I����V��^�E��e�w�u�u�w��F��I����W��^�E��e�d�e�e�g�l�F���Y���D��_�D��d�e�e�d�g�m�G��I����V��L����u�d�d�d�f�m�F��H����W��^�D��e�e�e�y�]�}�W��H����W��^�D��e�e�e�d�f�m�F��H���F�_�D��d�e�d�e�g�l�G��I����W��_�W���u�u�w�d�f�m�F��I����V��^�E��e�e�d�e�u�}�W���[����V��_�D��d�e�d�e�g�l�F��I����FǻN��D��d�e�e�e�g�l�G��I����W��^�D��y�_�u�u�f�l�F��H����V��_�E��d�e�d�e�f�l�[�ԜY���W��^�E��d�d�e�e�g�m�F��H����W�d��U���d�d�e�e�g�m�F��H����V��_�D��e�w�u�u�w��F��I����W��^�E��e�e�e�e�f�l�F���Y���D��_�E��d�e�d�e�f�m�G��I����W��L����u�d�d�d�g�m�G��I����V��^�E��d�d�e�y�]�}�W��H����W��_�E��e�e�e�d�g�m�G��I���F�_�D��d�d�e�d�g�l�G��I����V��_�W���u�u�w�d�f�l�F��I����W��^�E��d�d�d�d�u�}�W���[����W��^�D��d�e�d�e�g�l�F��I����FǻN��D��e�d�e�d�f�l�G��I����W��^�D��y�_�u�u�f�l�G��I����W��_�E��e�d�e�e�f�l�[�ԜY���W��_�D��e�d�e�d�g�m�G��I����V�d��U���d�d�d�d�g�m�F��H����V��^�D��e�w�u�u�w��F��H����W��^�E��e�e�d�e�g�l�F���Y���D��_�D��e�d�d�e�g�m�G��I����V��L����u�d�d�e�f�m�G��H����V��^�D��e�d�e�y�]�}�W��H����W��_�E��d�e�e�e�f�m�F��H���F�_�D��e�d�d�e�f�m�G��I����W��^�W���u�u�w�d�f�l�G��I����V��^�E��d�e�d�d�u�}�W���[����W��_�D��d�e�e�e�g�m�G��I����FǻN��D��e�d�d�d�f�m�G��I����V��^�E��y�_�u�u�f�l�G��H����W��_�D��d�d�e�d�f�m�[�ԜY���W��_�D��d�d�d�e�f�l�F��H����V�d��U���d�d�d�e�f�l�F��H����W��_�D��d�w�u�u�w��F��H����W��_�E��d�d�d�d�f�m�F���Y���D��_�D��e�d�d�e�f�m�F��H����W��L����u�d�d�e�f�m�G��H����V��_�E��d�d�e�y�]�}�W��H����V��^�D��e�d�d�d�g�m�F��H���F�_�D��d�e�d�e�g�l�F��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��d�e�d�d�u�}�W���[����W��_�E��e�e�d�d�f�m�G��H����FǻN��D��e�d�e�d�f�l�G��H����V��^�E��y�_�u�u�f�l�G��H����W��^�D��d�e�d�e�g�l�[�ԜY���W��_�E��d�d�d�d�f�l�F��I����W�d��U���d�d�d�d�f�m�F��I����W��^�E��d�w�u�u�w��F��H����V��^�D��d�d�e�e�g�m�F���Y���D��_�E��e�d�e�d�g�m�F��H����W��L����u�d�d�d�g�m�F��I����V��_�D��e�e�e�y�]�}�W��H����V��^�D��e�d�d�e�f�l�G��I���F�_�D��e�d�d�e�f�l�G��H����V��_�W���u�u�w�d�f�m�G��I����W��_�D��e�e�e�e�u�}�W���[����V��_�D��d�d�d�d�f�l�F��I����FǻN��D��d�e�d�d�g�l�F��I����W��_�E��y�_�u�u�f�l�F��I����W��_�D��e�e�d�d�f�m�[�ԜY���W��^�D��e�d�e�d�f�l�G��H����V�d��U���d�d�e�d�g�m�G��I����W��^�D��e�w�u�u�w��F��I����W��^�D��d�d�e�d�f�m�F���Y���D��_�E��d�e�d�e�g�l�F��I����V��L����u�d�d�d�f�m�G��I����W��_�D��e�d�e�y�]�}�W��H����V��_�E��e�d�d�e�f�m�G��I���F�_�D��e�d�d�d�f�l�G��H����W��^�W���u�u�w�d�f�m�G��H����V��_�D��e�e�d�d�u�}�W���[����V��_�D��d�d�d�d�f�m�G��H����FǻN��D��d�d�e�d�g�m�G��I����V��^�E��y�_�u�u�f�l�F��I����V��^�D��e�e�d�d�g�m�[�ԜY���W��_�E��e�e�e�e�f�l�G��H����W�d��U���d�d�e�d�f�m�G��I����W��^�E��d�w�u�u�w��F��H����V��_�E��d�d�e�d�f�l�F���Y���D��_�E��e�e�e�d�g�l�F��I����W��L����u�d�d�d�g�m�F��H����W��_�E��d�d�e�y�]�}�W��H����W��^�D��e�d�d�e�g�m�G��H���F�_�D��e�d�d�e�f�m�G��H����V��_�W���u�u�w�d�f�l�F��I����V��_�D��e�d�d�e�u�}�W���[����W��_�D��d�e�d�d�f�m�G��I����FǻN��D��d�e�d�d�f�m�G��H����V��_�E��y�_�u�u�f�l�F��H����V��^�D��e�e�d�e�f�l�[�ԜY���W��_�E��e�d�e�d�f�l�G��H����V�d��U���d�d�d�e�f�l�F��H����W��^�D��e�w�u�u�w��F��H����W��^�E��d�d�e�e�f�m�G���Y���D��_�D��e�e�d�d�f�m�F��I����V��L����u�d�d�d�f�m�G��H����V��_�E��d�d�e�y�]�}�W��H����V��_�E��e�d�d�e�g�m�G��H���F�_�D��d�e�e�e�g�m�G��H����V��_�W���u�u�w�d�f�l�F��I����W��_�D��d�e�d�d�u�}�W���[����V��^�E��e�e�e�d�f�m�F��H����FǻN��E��e�e�e�d�f�l�G��H����V��_�E��y�_�u�u�g�m�G��I����W��_�D��e�e�d�e�g�l�[�ԜY���V��^�E��d�e�d�d�f�l�G��H����V�d��U���e�e�e�e�f�m�F��H����W��^�D��d�w�u�u�w��G��I����W��_�E��d�d�e�e�g�l�G���Y���D��^�E��e�e�e�e�g�m�F��I����V��L����u�e�e�e�g�l�G��H����W��_�D��d�e�d�y�]�}�W��I����W��_�D��e�d�d�e�f�l�F��I���F�^�E��d�d�d�e�f�l�F��H����W��^�W���u�u�w�e�g�m�G��I����W��_�D��d�e�e�e�u�}�W���[����V��_�D��d�d�e�d�f�m�F��I����FǻN��E��e�d�d�e�f�l�G��H����V��^�E��y�_�u�u�g�m�G��H����W��^�D��e�d�d�d�g�l�[�ԜY���V��_�D��e�d�e�e�f�l�G��I����V�d��U���e�e�e�d�g�l�G��H����W��^�D��d�w�u�u�w��G��I����V��^�E��d�d�d�e�f�m�G���Y���D��^�D��d�e�d�e�g�m�F��H����V��L����u�e�e�e�f�l�G��I����W��_�E��e�d�d�y�]�}�W��I����W��^�D��d�d�d�e�g�l�F��I���F�^�E��d�d�e�d�f�l�G��H����V��^�W���u�u�w�e�g�l�G��H����W��_�D��e�d�d�e�u�}�W���[����W��^�D��d�e�d�d�f�l�G��H����FǻN��E��e�e�e�e�f�m�G��I����W��^�D��y�_�u�u�g�m�G��I����W��_�D��e�d�e�d�g�m�[�ԜY���V��^�E��e�e�d�e�f�l�G��H����V�d��U���e�e�d�e�f�m�G��H����W��^�E��d�w�u�u�w��G��H����W��^�D��d�d�e�e�f�l�F���Y���D��^�E��d�d�d�e�g�m�F��I����W��L����u�e�e�e�g�m�G��H����W��_�E��d�d�d�y�]�}�W��I����V��_�D��d�d�d�d�g�l�F��I���F�^�E��d�d�e�d�f�m�G��H����V��^�W���u�u�w�e�g�l�F��H����W��_�D��e�d�e�d�u�}�W���[����W��_�E��d�e�e�d�f�m�G��I����FǻN��E��e�e�d�e�g�l�G��I����V��^�D��y�_�u�u�g�m�G��H����W��^�D��d�d�d�e�g�l�[�ԜY���V��^�E��d�d�d�d�f�l�F��H����W�d��U���e�e�d�d�g�l�F��I����W��^�D��d�w�u�u�w��G��H����V��_�E��d�d�d�e�f�m�G���Y���D��^�E��e�d�d�d�f�l�F��H����V��L����u�e�e�e�g�l�G��I����W��_�E��e�d�e�y�]�}�W��I����W��^�E��d�d�d�d�g�l�F��I���F�^�E��d�d�e�d�f�m�G��H����V��^�W���u�u�w�e�g�l�F��I����V��_�D��e�e�d�e�u�}�W���[����W��_�E��e�e�e�d�f�l�F��H����FǻN��E��e�e�d�d�g�l�G��I����W��^�E��y�_�u�u�g�m�G��H����W��_�D��d�d�d�d�g�m�[�ԜY���V��^�D��e�d�e�e�g�m�G��I����V�d��U���e�e�d�d�f�m�F��I����V��^�E��d�w�u�u�w��G��H����V��^�D��e�e�e�d�g�m�F���Y���D��^�E��d�e�e�e�f�m�G��I����V��L����u�e�e�e�g�l�G��H����W��^�E��e�e�d�y�]�}�W��I����W��^�D��d�e�e�e�f�m�G��H���F�^�E��d�d�e�e�f�l�F��I����V��_�W���u�u�w�e�g�l�F��I����V��^�E��e�d�d�d�u�}�W���[����W��^�E��d�d�d�e�g�m�F��I����FǻN��E��e�e�d�d�g�m�F��I����V��^�E��y�_�u�u�g�m�G��H����W��^�E��e�d�d�e�f�m�[�ԜY���V��^�E��d�d�d�e�g�m�G��I����W�d��U���e�e�d�d�f�l�G��H����V��^�D��d�w�u�u�w��G��H����V��^�E��e�e�d�e�f�m�F���Y���D��^�E��e�d�e�e�f�m�G��H����W��L����u�e�e�e�g�m�F��H����W��^�E��d�e�d�y�]�}�W��I����V��^�E��e�e�e�e�g�l�F��I���F�^�E��d�e�e�e�g�m�G��I����W��_�W���u�u�w�e�g�l�G��I����V��^�E��e�e�d�d�u�}�W���[����W��_�E��e�d�e�e�g�l�G��I����FǻN��E��e�e�d�d�f�l�G��H����W��_�E��y�_�u�u�g�m�G��H����W��_�E��e�d�e�e�g�l�[�ԜY���V��^�E��e�d�e�e�g�m�G��I����W�d��U���e�e�d�e�f�m�G��H����V��_�D��e�w�u�u�w��G��H����V��^�E��e�e�d�d�g�l�G���Y���D��^�E��d�e�e�d�f�l�G��H����V��L����u�e�e�e�g�m�G��I����V��^�E��e�d�d�y�]�}�W��I����W��^�D��d�e�e�d�g�m�G��H���F�^�E��d�d�e�e�f�l�F��I����V��_�W���u�u�w�e�g�m�F��H����W��^�E��e�e�e�d�u�}�W���[����V��_�D��d�d�d�e�g�m�G��I����FǻN��E��e�d�e�e�g�l�F��H����V��_�E��y�_�u�u�g�m�G��I����W��^�E��d�e�e�e�g�l�[�ԜY���V��_�E��d�e�e�d�g�m�F��I����V�d��U���e�e�e�e�f�m�G��H����V��^�D��d�w�u�u�w��G��I����V��_�E��e�e�e�d�f�l�G���Y���D��^�D��e�d�e�e�f�m�G��I����V��L����u�e�e�e�f�m�F��H����W��^�E��d�e�d�y�]�}�W��I����V��^�E��e�e�e�d�g�l�F��H���F�^�E��e�e�e�e�g�l�G��I����W��^�W���u�u�w�e�g�m�G��I����V��^�E��d�d�d�d�u�}�W���[����V��_�D��e�e�e�e�g�m�F��I����FǻN��E��e�e�d�d�g�l�G��I����V��_�D��y�_�u�u�g�m�G��H����W��_�E��d�e�d�d�g�l�[�ԜY���V��^�D��e�e�d�e�g�m�F��H����W�d��U���e�e�e�d�g�l�G��H����V��^�D��d�w�u�u�w��G��I����W��_�E��e�e�e�d�f�l�F���Y���D��^�E��d�d�d�e�g�m�G��I����W��L����u�e�e�e�g�l�G��H����V��^�E��d�d�e�y�]�}�W��I����W��_�E��d�e�e�d�g�l�F��I���F�^�E��e�d�d�d�g�m�F��I����W��_�W���u�u�w�e�g�m�G��I����V��^�E��d�d�e�e�u�}�W���[����V��^�E��d�d�e�e�g�m�F��H����FǻN��E��e�e�e�e�g�m�G��I����V��^�D��y�_�u�u�f�l�F��H����V��_�E��d�e�d�e�g�m�[�ԜY���W��_�E��e�d�d�e�g�m�F��I����V�d��U���d�d�d�d�g�m�F��I����V��^�D��d�w�u�u�w��F��H����V��_�E��e�e�e�d�f�m�G���Y���D��_�D��e�e�e�e�f�l�G��I����V��L����u�d�d�d�f�m�F��I����V��^�E��e�d�d�y�]�}�W��H����W��_�E��e�e�e�d�g�l�F��I���F�_�D��e�d�d�e�f�m�G��I����W��^�W���u�u�w�d�f�l�G��H����V��^�E��e�e�e�e�u�}�W���[����W��^�E��e�d�d�e�g�m�G��H����FǻN��D��d�d�e�d�g�l�F��I����V��_�D��y�_�u�u�f�l�F��I����W��_�E��d�e�e�d�g�m�[�ԜY���W��_�E��e�d�e�e�g�m�G��H����W�d��U���d�d�d�e�g�l�F��H����V��_�D��e�w�u�u�w��F��H����W��^�E��e�e�d�d�g�l�G���Y���D��_�E��e�d�e�e�f�l�G��H����V��L����u�d�d�d�g�l�F��H����W��^�D��d�e�d�y�]�}�W��H����W��_�D��d�e�e�e�f�l�F��H���F�_�D��d�e�e�d�g�m�F��I����W��_�W���u�u�w�d�f�l�F��I����W��^�E��e�e�d�e�u�}�W���[����W��_�E��d�d�e�e�g�l�G��H����FǻN��D��d�e�e�d�f�m�G��H����W��^�D��y�_�u�u�f�l�F��I����V��_�E��e�e�d�d�g�m�[�ԜY���W��^�E��e�e�d�d�g�m�G��H����V�d��U���d�d�d�e�f�l�F��I����V��^�D��e�w�u�u�w��F��H����W��_�D��e�e�d�d�g�m�F���Y���D��_�E��e�d�e�e�f�m�G��H����V��L����u�d�d�d�g�l�F��I����W��^�E��d�e�e�y�]�}�W��H����W��^�D��d�e�e�e�g�m�F��I���F�_�D��e�e�d�d�g�l�F��I����V��^�W���u�u�w�d�f�l�G��I����W��^�E��d�d�e�d�u�}�W���[����W��_�D��d�e�e�e�g�m�F��I����FǻN��D��d�e�e�d�f�l�F��H����V��_�D��y�_�u�u�f�l�F��I����W��^�E��e�d�e�d�f�m�[�ԜY���W��^�D��e�e�e�e�g�m�G��H����W�d��U���d�d�d�e�f�m�G��I����V��_�E��d�w�u�u�w��F��H����W��^�E��e�e�e�e�f�m�G���Y���D��_�E��d�e�d�e�f�m�G��I����W��L����u�d�d�d�g�m�F��H����W��^�E��e�d�e�y�]�}�W��H����V��_�E��d�e�e�e�g�l�G��I���F�_�D��e�e�e�e�f�m�G��I����V��^�W���u�u�w�d�f�l�G��H����V��^�E��d�e�d�d�u�}�W���[����W��^�D��e�d�e�e�g�m�G��H����FǻN��D��d�e�e�e�f�m�G��I����V��^�E��y�_�u�u�f�l�F��I����W��_�E��e�e�e�e�f�l�[�ԜY���W��^�E��d�d�d�e�g�m�G��I����W�d��U���d�d�d�e�g�l�G��I����W��_�D��d�w�u�u�w��F��H����W��^�E��d�d�d�d�g�m�F���Y���D��_�E��e�d�e�e�g�l�F��H����V��L����u�d�d�d�g�m�F��I����W��_�D��e�e�e�y�]�}�W��H����V��^�D��d�d�d�d�f�l�G��H���F�_�D��e�e�e�e�f�m�F��H����W��^�W���u�u�w�d�f�l�G��H����W��_�D��e�d�d�e�u�}�W���[����W��^�D��e�e�d�d�f�l�G��I����FǻN��D��d�e�e�e�g�m�F��I����W��_�E��y�_�u�u�f�l�F��I����W��^�D��d�e�d�d�f�m�[�ԜY���W��^�D��d�d�d�e�f�l�F��I����V�d��U���d�d�d�e�f�m�G��H����W��^�E��d�w�u�u�w��F��H����V��^�D��d�d�d�d�g�m�G���Y���D��_�E��d�d�e�d�g�l�F��H����W��L����u�d�d�d�g�l�G��H����W��_�E��d�e�e�y�]�}�W��H����W��^�E��d�d�d�d�g�m�F��I���F�_�D��e�e�e�e�f�m�G��H����V��_�W���u�u�w�d�f�l�G��H����W��_�D��e�e�d�e�u�}�W���[����W��_�E��d�e�d�d�f�m�F��I����FǻN��D��d�e�d�e�g�m�G��I����V��^�E��y�_�u�u�f�l�F��H����W��^�D��d�d�d�e�f�m�[�ԜY���W��^�D��e�d�d�e�f�l�F��I����W�d��U���d�d�d�d�g�m�F��H����W��_�E��e�w�u�u�w��F��H����V��^�E��d�d�e�d�g�l�F���Y���D��_�E��d�e�e�e�g�m�F��I����W��L����u�d�d�d�g�m�G��I����W��_�D��e�d�d�y�]�}�W��H����V��_�E��e�d�d�d�f�l�F��I���F�_�D��d�d�d�d�g�m�F��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��e�d�e�d�u�}�W���[����W��^�E��e�d�d�d�f�m�G��H����FǻN��D��d�e�d�d�f�m�G��H����V��^�D��y�_�u�u�f�l�F��H����W��^�D��d�d�e�d�g�m�[�ԜY���W��^�D��d�d�e�d�f�l�F��I����V�d��U���d�d�d�d�f�l�F��H����W��^�D��e�w�u�u�w��F��H����W��^�D��d�d�e�d�f�m�G���Y���D��_�D��d�e�e�e�f�l�F��I����V��L����u�d�d�d�f�m�G��H����V��_�E��d�d�d�y�]�}�W��H����V��^�D��e�d�d�d�g�l�F��I���F�_�D��e�d�d�d�g�l�F��H����W��^�W���u�u�w�d�f�l�G��H����V��_�D��d�e�d�e�u�}�W���[����W��^�E��e�e�d�d�f�m�F��H����FǻN��D��d�d�d�e�f�l�G��I����V��^�D��y�_�u�u�f�l�F��H����V��_�D��d�e�d�e�g�l�[�ԜY���W��_�D��d�e�e�d�f�l�F��I����W�d��U���d�d�d�d�g�l�G��H����W��^�D��d�w�u�u�w��F��H����W��^�E��d�d�e�d�f�l�F���Y���D��_�D��e�d�e�e�f�l�F��I����W��L����u�d�d�d�f�m�F��H����W��_�E��e�e�e�y�]�}�W��H����W��^�E��d�d�d�d�g�l�G��I���F�_�D��d�e�d�e�g�m�G��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�e�d�e�u�}�W���[����W��_�D��e�d�d�d�f�m�F��H����FǻN��D��d�d�d�d�g�l�F��I����V��^�D��y�_�u�u�g�m�G��I����V��^�D��d�e�d�d�g�m�[�ԜY���V��^�E��e�e�d�d�f�l�F��H����W�d��U���e�e�e�e�g�l�G��I����W��^�D��e�w�u�u�w��G��I����V��^�D��d�d�e�d�f�m�G���Y���D��^�E��d�e�d�e�g�l�F��I����W��L����u�e�e�e�g�m�F��H����V��_�D��e�d�e�y�]�}�W��I����W��^�D��e�d�d�d�f�m�G��H���F�^�E��e�e�e�e�g�l�G��H����V��^�W���u�u�w�e�g�m�G��H����V��_�D��e�d�e�d�u�}�W���[����V��_�E��e�d�e�d�f�m�G��I����FǻN��E��e�e�d�d�f�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��_�D��d�d�d�e�f�m�[�ԜY���V��^�E��d�e�d�d�f�l�F��H����V�d��U���e�e�e�d�g�m�G��I����W��_�D��d�w�u�u�w��G��I����W��_�D��d�d�e�e�f�l�F���Y���D��^�E��e�e�d�e�g�l�F��I����W��L����u�e�e�e�g�m�F��H����V��_�D��d�e�d�y�]�}�W��I����V��_�D��e�d�d�d�f�m�G��I���F�^�E��d�e�e�e�f�m�F��H����V��_�W���u�u�w�e�g�m�F��H����W��_�D��d�e�d�d�u�}�W���[����V��^�D��d�d�d�d�f�m�F��I����FǻN��E��e�e�d�d�f�l�G��H����V��_�D��y�_�u�u�g�m�G��H����V��_�D��d�e�e�e�f�l�[�ԜY���V��^�D��d�d�e�d�f�l�F��I����V�d��U���e�e�e�d�f�m�G��I����W��^�D��d�w�u�u�w��G��I����W��_�E��d�d�d�e�g�m�F���Y���D��^�D��e�e�d�d�f�l�F��H����V��L����u�e�e�e�f�m�G��H����W��_�E��e�e�e�y�]�}�W��I����V��_�D��e�d�d�d�g�l�F��H���F�^�E��e�e�e�e�f�m�G��H����V��_�W���u�u�w�e�g�m�G��H����V��_�D��d�d�d�e�u�}�W���[����V��^�D��d�e�e�d�f�l�F��H����FǻN��E��e�d�e�e�f�m�G��I����W��^�D��y�_�u�u�g�m�G��I����V��^�D��d�e�d�e�g�l�[�ԜY���V��_�D��e�d�d�e�f�l�F��H����W�d��U���e�e�e�e�f�m�G��H����W��_�E��e�w�u�u�w��G��I����V��_�D��d�d�d�e�f�l�F���Y���D��^�D��d�d�e�d�f�m�F��H����V��L����u�e�e�e�f�m�F��H����V��_�D��d�d�e�y�]�}�W��I����V��^�D��e�d�d�d�f�l�G��H���F�^�E��e�d�d�e�f�l�G��H����V��^�W���u�u�w�e�g�m�G��H����V��_�D��d�e�e�d�u�}�W���[����V��^�E��d�e�d�d�f�l�F��H����FǻN��E��e�d�d�e�g�l�F��H����W��^�E��y�_�u�u�g�m�G��H����V��^�D��d�d�d�d�f�l�[�ԜY���V��_�E��d�d�e�e�f�l�F��H����V�d��U���e�e�e�e�g�m�F��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�m�F���Y���D��^�D��e�e�d�d�g�l�G��I����W��L����u�e�e�e�f�l�G��I����W��^�E��d�d�d�y�]�}�W��I����V��_�D��d�e�e�e�g�l�F��H���F�^�E��e�d�d�e�f�l�G��I����W��_�W���u�u�w�e�g�m�G��H����V��^�E��e�d�d�d�u�}�W���[����V��_�E��d�d�e�e�g�m�F��H����FǻN��E��e�d�e�d�f�l�F��I����V��_�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�d�g�l�[�ԜY���V��_�D��e�e�d�e�g�m�G��H����W�d��U���e�e�e�e�f�l�F��I����V��^�E��d�w�u�u�w��G��I����W��^�D��e�e�e�d�f�l�G���Y���D��^�D��e�d�e�e�g�m�G��I����W��L����u�e�e�e�f�m�G��I����V��^�D��e�e�e�y�]�}�W��I����V��_�D��e�e�e�e�f�m�F��H���F�^�E��e�e�d�e�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�d�d�d�u�}�W���[����V��^�D��d�e�e�e�g�m�G��H����FǻN��E��e�d�e�e�g�l�F��H����V��^�D��y�_�u�u�g�m�G��I����V��_�E��e�d�d�e�f�l�[�ԜY���V��^�D��d�d�e�e�g�m�G��H����W�d��U���e�e�e�d�f�l�G��I����V��_�E��e�w�u�u�w��G��I����V��^�D��e�e�e�d�g�l�G���Y���D��^�E��e�e�d�d�f�m�G��I����W��L����u�e�e�e�g�l�G��H����V��^�D��e�d�e�y�]�}�W��I����W��_�D��d�e�e�e�f�m�G��H���F�^�E��d�e�e�d�f�m�G��I����V��^�W���u�u�w�e�g�m�F��I����W��^�E��d�e�e�d�u�}�W���[����V��^�E��e�e�d�e�g�m�F��H����FǻN��E��e�e�d�e�g�m�G��I����V��^�D��y�_�u�u�g�m�G��I����V��_�E��e�d�d�d�f�l�[�ԜY���V��^�D��d�e�d�d�g�m�G��H����W�d��U���e�e�e�d�f�l�F��H����V��_�D��e�w�u�u�w��G��I����V��_�E��e�e�e�d�f�m�F���Y���D��^�E��d�e�d�d�g�l�G��I����W��L����u�e�e�e�g�m�F��H����W��^�D��d�d�e�y�]�}�W��I����V��^�D��d�e�e�e�g�m�G��H���F�^�E��d�e�e�d�f�l�G��I����V��_�W���u�u�w�e�g�m�G��H����V��^�E��e�e�d�d�u�}�W���[����V��_�E��d�e�d�e�g�l�G��H����FǻN��E��e�e�d�e�g�l�G��H����W��^�E��y�_�u�u�g�m�G��H����V��^�E��e�e�e�d�g�m�[�ԜY���V��^�E��d�e�d�e�g�m�G��I����V�d��U���e�e�e�e�g�m�F��H����V��^�E��e�w�u�u�w��G��I����W��_�D��e�e�d�e�g�m�G���Y���D��^�E��e�e�d�d�f�l�G��H����V��L����u�e�e�e�g�m�F��H����W��^�E��d�d�e�y�]�}�W��I����V��^�D��e�e�e�e�g�m�F��H���F�^�E��e�d�d�e�f�m�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�d�u�}�W���[����V��^�E��e�d�d�e�g�l�G��H����FǻN��E��e�e�e�d�g�m�G��H����W��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�f�l�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�G��I����V��_�D��d�w�u�u�w��F��H����V��^�D��e�e�e�d�f�m�F���Y���D��_�D��e�e�e�d�f�m�G��I����V��L����u�d�d�d�f�l�G��I����V��^�D��e�e�e�y�]�}�W��H����W��^�E��e�e�e�e�f�l�G��I���F�_�D��d�e�e�e�f�m�G��I����W��_�W���u�u�w�d�f�l�F��H����W��^�E��d�e�e�e�u�}�W���[����W��^�E��d�e�e�e�g�m�F��H����FǻN��D��d�d�e�d�f�m�G��H����V��^�D��y�_�u�u�f�l�F��I����W��^�E��e�d�e�d�f�m�[�ԜY���W��_�D��d�e�d�d�g�m�G��I����W�d��U���d�d�d�d�f�m�F��I����V��_�D��d�w�u�u�w��F��H����V��^�D��e�e�e�d�f�m�G���Y���D��_�D��d�e�e�d�f�m�G��I����V��L����u�d�d�d�f�m�F��I����V��^�D��e�d�e�y�]�}�W��H����V��_�D��e�e�e�e�f�m�G��H���F�_�D��d�e�d�e�f�l�F��I����W��_�W���u�u�w�d�f�l�F��I����V��^�E��e�d�d�d�u�}�W���[����W��_�D��d�e�e�e�g�m�G��H����FǻN��D��d�d�d�d�g�m�F��I����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�d�d�e�f�l�[�ԜY���W��_�D��d�e�d�e�g�m�G��I����W�d��U���d�d�d�e�f�l�G��H����V��_�D��d�w�u�u�w��F��H����V��^�E��e�e�e�e�f�m�F���Y���D��_�D��e�e�e�d�f�l�G��I����V��L����u�d�d�d�f�l�F��I����W��^�D��e�e�e�y�]�}�W��H����W��^�D��d�e�e�e�g�l�F��H���F�_�D��e�e�e�e�g�m�G��I����W��_�W���u�u�w�d�f�l�G��I����V��^�E��d�d�e�e�u�}�W���[����W��^�D��d�e�e�e�g�m�F��I����FǻN��D��d�d�d�e�g�l�G��I����V��^�D��y�_�u�u�f�l�F��H����V��^�E��e�e�e�d�g�m�[�ԜY���W��_�E��e�d�e�d�g�m�G��I����W�d��U���d�d�d�e�g�m�F��H����V��^�E��e�w�u�u�w��F��H����V��_�E��e�e�e�d�g�l�F���Y���D��_�D��d�d�e�d�g�m�G��I����V��L����u�d�d�d�f�m�F��H����V��^�E��d�d�e�y�]�}�W��H����V��^�D��e�e�e�e�g�l�G��I���F�_�D��e�d�d�d�g�l�G��I����W��^�W���u�u�w�d�f�l�G��H����W��^�E��e�e�d�d�u�}�W���[����W��_�E��e�e�d�e�g�m�G��H����FǻN��D��d�d�e�d�f�l�F��H����V��_�D��y�_�u�u�f�l�F��I����V��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�d�d�g�m�G��I����W�d��U���d�d�d�e�f�m�F��I����V��^�E��d�w�u�u�w��F��H����V��^�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�e�e�f�m�F��H����W��L����u�d�d�d�f�m�F��H����W��_�D��e�e�e�y�]�}�W��H����V��_�D��d�d�d�d�f�l�F��I���F�_�D��e�d�d�e�f�m�G��H����W��_�W���u�u�w�d�f�l�G��H����V��_�D��d�d�d�d�u�}�W���[����W��_�E��e�d�e�d�f�l�F��H����FǻN��D��d�d�e�d�f�m�G��I����W��_�E��y�_�u�u�f�l�F��I����V��_�D��d�d�e�d�f�l�[�ԜY���W��_�E��e�e�e�e�f�l�F��I����V�d��U���d�d�d�e�g�m�F��I����W��_�E��e�w�u�u�w��F��H����V��^�E��d�d�d�e�f�m�G���Y���D��_�D��e�d�e�e�g�l�F��H����W��L����u�d�d�d�f�l�G��H����W��_�D��e�e�e�y�]�}�W��H����W��^�D��d�d�d�d�f�l�F��I���F�_�D��e�e�d�d�g�l�F��H����W��_�W���u�u�w�d�f�l�G��I����W��_�D��e�e�e�d�u�}�W���[����W��^�D��e�d�d�d�f�l�G��H����FǻN��D��d�d�d�d�f�l�F��H����W��_�D��y�_�u�u�f�l�F��H����W��_�D��d�d�e�e�f�l�[�ԜY���W��_�E��d�d�e�e�f�l�F��I����V�d��U���d�d�d�e�f�m�F��H����W��_�E��d�w�u�u�w��F��H����V��^�D��d�d�d�e�g�l�F���Y���D��_�D��e�e�e�e�f�m�F��H����V��L����u�d�d�d�f�l�G��I����V��_�E��d�d�d�y�]�}�W��H����W��^�E��d�d�d�d�g�l�F��I���F�_�D��e�d�e�d�g�l�G��H����W��^�W���u�u�w�d�f�l�G��H����V��_�D��d�d�d�e�u�}�W���[����W��_�D��e�e�e�d�f�l�F��I����FǻN��D��d�d�e�e�g�l�G��I����W��_�E��y�_�u�u�f�l�F��I����V��_�D��d�e�d�d�g�l�[�ԜY���W��_�E��e�d�d�e�f�l�F��H����V�d��U���d�d�d�d�g�m�G��I����W��^�E��d�w�u�u�w��F��H����V��^�E��d�d�d�d�g�l�F���Y���D��_�D��d�e�d�e�f�m�F��H����W��L����u�d�d�d�f�m�G��I����V��_�E��e�d�d�y�]�}�W��H����V��_�E��e�d�d�d�g�l�G��I���F�_�D��d�d�d�d�g�m�F��H����W��^�W���u�u�w�d�f�l�F��H����V��_�D��d�d�d�d�u�}�W���[����W��_�D��e�e�e�d�f�l�F��H����FǻN��D��d�d�e�d�g�l�G��H����W��_�E��y�_�u�u�f�l�F��I����V��^�D��d�e�e�d�g�m�[�ԜY���W��_�E��d�e�d�d�f�l�F��I����W�d��U���d�d�d�d�g�l�G��I����W��^�D��e�w�u�u�w��F��H����W��_�E��d�d�d�d�f�l�G���Y���D��_�D��d�e�e�d�g�m�F��H����W��L����u�d�d�d�f�l�F��H����V��_�E��d�e�e�y�]�}�W��H����W��_�E��e�d�d�d�g�m�F��H���F�_�D��d�d�e�d�g�m�F��H����V��^�W���u�u�w�d�f�l�F��I����W��_�D��d�d�d�e�u�}�W���[����W��_�D��e�d�d�d�f�l�F��H����FǻN��D��d�d�d�d�g�l�G��I����W��_�D��y�_�u�u�f�l�F��H����V��_�D��d�e�d�e�g�m�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����V�d��U���e�e�e�e�g�m�G��I����W��^�E��d�w�u�u�w��G��I����V��_�D��d�d�d�d�g�l�F���Y���D��^�E��e�e�d�e�f�l�F��H����W��L����u�e�e�e�g�m�G��I����W��_�E��d�e�e�y�]�}�W��I����V��^�D��d�d�d�d�g�l�F��I���F�^�E��e�e�e�d�f�m�G��H����W��^�W���u�u�w�e�g�m�G��H����V��_�D��d�e�d�d�u�}�W���[����V��_�E��e�e�d�d�f�l�F��I����FǻN��E��e�e�e�e�f�m�F��I����W��_�E��y�_�u�u�g�m�G��I����W��_�D��d�e�d�e�f�m�[�ԜY���V��^�D��e�e�d�e�f�l�F��H����V�d��U���e�e�e�e�f�m�G��H����W��^�D��e�w�u�u�w��G��I����V��_�E��d�d�d�d�f�l�F���Y���D��^�E��d�e�d�d�g�m�F��H����V��L����u�e�e�e�g�m�F��H����V��_�D��e�d�e�y�]�}�W��I����W��^�D��e�d�d�d�f�m�F��I���F�^�E��e�e�e�e�f�m�F��H����V��^�W���u�u�w�e�g�m�G��H����V��_�D��e�d�e�e�u�}�W���[����V��^�E��d�d�e�d�f�l�G��I����FǻN��E��e�e�d�e�f�m�G��I����W��_�D��y�_�u�u�g�m�G��H����W��^�D��d�d�e�d�f�l�[�ԜY���V��^�E��e�d�d�e�f�l�F��I����W�d��U���e�e�e�e�g�m�F��I����W��_�E��e�w�u�u�w��G��I����W��_�E��d�d�d�e�g�l�G���Y���D��^�E��d�d�d�d�f�l�F��H����V��L����u�e�e�e�g�l�F��H����W��_�D��d�d�e�y�]�}�W��I����W��^�E��d�d�d�d�f�l�G��I���F�^�E��e�d�e�e�f�l�F��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��e�d�e�e�u�}�W���[����V��_�E��d�e�d�d�f�l�G��H����FǻN��E��e�e�d�e�g�m�F��H����W��^�D��y�_�u�u�g�m�G��H����V��^�D��d�d�e�e�f�l�[�ԜY���V��^�D��d�e�e�e�f�l�F��I����W�d��U���e�e�e�e�f�l�F��I����W��_�E��e�w�u�u�w��G��I����V��^�E��d�d�d�d�f�m�F���Y���D��^�E��d�e�e�e�f�m�F��H����W��L����u�e�e�e�g�l�F��H����V��_�D��d�d�e�y�]�}�W��I����W��_�D��d�d�d�d�f�m�F��H���F�^�E��e�d�e�e�f�l�G��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�e�d�d�u�}�W���[����V��_�D��e�e�d�d�f�l�F��I����FǻN��E��e�e�d�d�f�l�G��I����W��_�E��y�_�u�u�g�m�G��H����W��^�D��d�d�d�e�g�m�[�ԜY���V��^�D��e�e�d�d�f�l�F��H����V�d��U���e�e�e�e�f�l�G��I����W��_�D��e�w�u�u�w��G��I����W��^�E��e�e�e�e�g�m�G���Y���D��^�E��d�e�e�e�g�l�G��I����W��L����u�e�e�e�g�l�F��H����V��^�E��e�d�d�y�]�}�W��I����W��_�D��e�e�e�e�g�m�F��H���F�^�E��e�d�e�d�g�m�F��I����V��_�W���u�u�w�e�g�m�G��I����V��^�E��e�d�e�d�u�}�W���[����V��_�D��d�e�d�e�g�m�G��H����FǻN��E��e�e�d�d�f�m�F��H����V��_�D��y�_�u�u�g�m�G��H����V��_�E��e�e�e�d�g�l�[�ԜY���V��^�D��d�e�e�e�g�m�G��H����V�d��U���e�e�e�e�f�m�G��H����V��^�E��e�w�u�u�w��G��I����V��_�E��e�e�e�e�g�m�G���Y���D��^�E��e�d�d�d�g�m�G��I����V��L����u�e�e�e�g�l�G��H����V��^�E��d�d�e�y�]�}�W��I����W��_�E��d�e�e�e�g�l�G��H���F�^�E��e�d�d�d�f�l�F��I����W��^�W���u�u�w�e�g�m�G��H����W��^�E��e�d�d�d�u�}�W���[����V��_�D��e�e�e�e�g�m�G��I����FǻN��E��e�e�d�e�f�l�G��H����V��_�E��y�_�u�u�g�m�G��H����W��^�E��e�e�d�d�f�l�[�ԜY���V��^�D��e�e�d�e�g�m�G��I����V�d��U���e�e�e�e�g�l�F��I����V��^�E��e�w�u�u�w��G��I����W��_�D��e�e�e�d�g�l�G���Y���D��^�E��d�e�e�e�f�m�G��I����V��L����u�e�e�e�g�l�F��I����V��^�E��d�d�e�y�]�}�W��I����W��_�D��e�e�e�e�g�m�F��I���F�^�E��e�e�e�d�g�m�F��I����V��_�W���u�u�w�e�g�m�G��I����V��^�E��d�d�e�d�u�}�W���[����V��^�D��e�d�d�e�g�m�F��I����FǻN��E��e�e�d�e�g�l�G��H����V��_�E��y�_�u�u�g�m�G��H����V��^�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�e�d�e�g�m�G��I����V�d��U���e�e�e�e�g�m�F��H����V��^�D��e�w�u�u�w��G��I����V��_�E��e�e�e�d�f�m�F���Y���D��^�E��d�d�d�d�g�l�G��I����V��L����u�e�e�e�g�m�F��I����W��^�E��d�e�e�y�]�}�W��I����V��^�E��d�e�e�e�g�m�F��H���F�^�E��e�d�e�e�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��d�d�d�e�u�}�W���[����V��_�D��e�d�d�e�g�m�F��H����FǻN��E��e�e�e�e�f�m�G��H����V��_�D��y�_�u�u�g�m�G��I����W��^�E��e�e�e�d�f�l�[�ԜY���V��^�D��d�e�e�e�g�m�G��H����V�d��U���e�e�e�e�f�m�F��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�d�g�m�G���Y���D��^�E��d�d�d�d�g�l�G��I����V��L����u�e�e�e�g�m�F��I����W��^�E��e�e�e�y�]�}�W��I����V��_�E��d�e�e�e�g�m�F��H���F�^�E��e�e�e�e�g�m�F��I����V��_�W���u�u�w�e�g�m�G��I����V��^�E��d�d�d�d�u�}�W���[����V��^�D��d�e�d�e�g�m�F��H����FǻN��E��e�e�e�e�g�l�F��I����V��_�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�d�g�m�[�ԜY���V��^�E��e�d�d�d�g�m�G��I����V�d��U���e�e�e�e�g�m�F��I����V��^�D��d�w�u�u�w��G��I����V��^�E��e�e�e�d�f�m�G���Y���D��_�D��d�d�d�e�f�l�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��d�e�e�y�]�}�W��H����W��_�D��d�e�e�e�g�m�G��I���F�_�D��d�d�e�e�g�m�G��I����V��^�W���u�u�w�d�f�l�F��I����W��^�E��d�d�d�e�u�}�W���[����W��_�D��d�d�d�e�g�m�F��I����FǻN��D��d�d�d�e�f�l�F��I����V��_�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��e�e�e�d�g�m�G��I����V�d��U���d�d�d�d�f�m�G��H����V��^�E��e�w�u�u�w��F��H����V��_�D��e�e�e�d�g�m�F���Y���D��_�D��e�e�d�d�f�l�G��I����V��L����u�d�d�d�f�l�F��H����W��^�E��e�d�e�y�]�}�W��H����W��_�D��e�e�e�e�g�m�G��I���F�_�D��d�e�d�d�f�m�F��I����V��_�W���u�u�w�d�f�l�F��H����V��^�E��d�e�e�d�u�}�W���[����W��^�D��d�d�d�e�g�m�G��H����FǻN��D��d�d�d�d�f�m�F��H����V��_�E��y�_�u�u�f�l�F��H����W��_�E��e�e�d�d�f�m�[�ԜY���W��_�E��e�e�e�d�g�m�G��H����V�d��U���d�d�d�d�g�l�F��I����V��^�D��e�w�u�u�w��F��H����W��_�D��e�e�e�e�f�l�G���Y���D��_�D��e�d�e�d�g�l�G��I����V��L����u�d�d�d�f�l�G��I����V��^�E��e�e�e�y�]�}�W��H����W��^�E��d�e�e�e�g�l�F��H���F�_�D��d�e�d�e�g�l�G��I����W��_�W���u�u�w�d�f�l�F��I����V��^�E��e�e�e�d�u�}�W���[����W��^�D��e�e�e�e�g�m�G��H����FǻN��D��d�d�d�e�f�m�G��H����V��^�E��y�_�u�u�f�l�F��H����W��_�E��e�e�d�e�g�l�[�ԜY���W��_�E��d�e�d�d�g�m�G��I����W�d��U���d�d�d�d�g�m�G��I����V��^�D��d�w�u�u�w��F��H����V��_�E��e�e�e�e�f�m�G���Y���D��_�D��e�e�e�e�g�m�G��I����V��L����u�d�d�d�f�m�F��H����W��^�E��e�e�d�y�]�}�W��H����V��_�D��d�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����W��^�E��e�e�d�e�u�}�W���[����W��_�D��d�d�e�e�g�m�G��H����FǻN��D��d�d�e�d�f�l�G��I����V��^�D��y�_�u�u�f�l�F��I����V��^�E��e�e�e�e�f�l�[�ԜY���W��_�D��e�d�d�e�g�m�G��I����W�d��U���d�d�d�d�f�l�G��I����V��^�E��d�w�u�u�w��F��H����W��_�E��e�e�e�e�g�m�F���Y���D��_�D��d�d�e�e�f�m�F��H����W��L����u�d�d�d�f�m�F��I����W��_�D��d�e�d�y�]�}�W��H����V��_�D��d�d�d�d�f�l�F��I���F�_�D��d�d�d�e�g�m�F��H����W��^�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�e�u�}�W���[����W��_�D��d�e�d�d�f�l�F��H����FǻN��D��d�d�e�d�f�m�G��H����W��_�D��y�_�u�u�f�l�F��I����V��_�D��d�d�d�e�g�m�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��H����W��_�E��e�w�u�u�w��F��H����V��_�D��d�d�d�d�g�m�G���Y���D��_�D��e�e�d�d�f�m�F��H����V��L����u�d�d�d�f�l�G��I����W��_�D��e�d�d�y�]�}�W��H����W��^�D��d�d�d�d�f�l�G��I���F�_�D��d�e�e�d�f�l�G��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��d�e�e�d�u�}�W���[����W��^�D��d�d�e�d�f�l�F��I����FǻN��D��d�d�d�e�f�m�F��H����W��_�D��y�_�u�u�f�l�F��H����W��_�D��d�d�e�d�g�m�[�ԜY���W��_�E��e�e�e�d�f�l�F��I����W�d��U���d�d�d�d�g�l�F��I����W��_�D��e�w�u�u�w��F��H����W��_�E��d�d�d�d�f�m�F���Y���D��_�D��e�d�e�d�g�l�F��H����V��L����u�d�d�d�f�l�G��I����V��_�D��e�d�d�y�]�}�W��H����W��_�E��e�d�d�d�f�m�G��H���F�_�D��d�e�e�e�f�m�G��H����V��^�W���u�u�w�d�f�l�F��I����W��_�D��d�d�e�d�u�}�W���[����W��^�E��e�d�d�d�f�l�F��I����FǻN��D��d�d�d�d�f�l�G��I����W��_�E��y�_�u�u�f�l�F��H����V��^�D��d�d�e�e�g�l�[�ԜY���W��_�E��e�e�e�e�f�l�F��I����V�d��U���d�d�d�d�g�l�G��I����W��_�E��d�w�u�u�w��F��H����W��^�D��d�d�d�d�g�l�G���Y���D��_�D��d�d�e�e�g�l�F��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�e�d�y�]�}�W��H����W��_�D��e�d�d�d�f�m�F��I���F�_�D��d�d�e�e�g�l�F��H����V��^�W���u�u�w�d�f�l�F��I����V��_�D��d�e�d�e�u�}�W���[����W��_�D��e�e�e�d�f�l�F��H����FǻN��D��d�d�d�e�f�m�F��H����W��^�D��y�_�u�u�f�l�F��H����W��^�D��d�d�e�d�f�l�[�ԜY���W��_�D��e�d�e�e�f�l�F��I����W�d��U���d�d�d�d�f�l�F��H����W��_�E��d�w�u�u�w��F��H����W��_�D��d�d�d�d�g�m�F���Y���D��_�D��e�d�e�e�g�m�F��H����V��L����u�d�d�d�f�l�F��I����W��_�D��d�d�d�y�]�}�W��H����W��^�D��d�d�d�d�f�m�F��H���F�_�D��d�d�e�d�g�l�F��H����V��^�W���u�u�w�d�f�l�F��I����V��_�D��d�e�d�e�u�}�W���[����W��_�D��e�e�e�d�f�l�F��H����FǻN��D��d�d�d�d�g�m�G��H����W��^�E��y�_�u�u�f�l�F��H����W��_�D��d�d�e�d�g�l�[�ԜY���W��_�D��d�e�d�e�f�l�F��I����W�d��U���d�d�d�d�f�l�G��H����W��_�E��e�w�u�u�w��F��H����W��^�D��d�d�d�d�g�l�F���Y���D��^�E��e�e�e�e�g�m�F��H����W��L����u�e�e�e�g�m�G��H����V��_�D��e�e�e�y�]�}�W��I����V��^�D��d�d�d�d�f�m�G��H���F�^�E��e�e�e�e�g�l�G��H����V��^�W���u�u�w�e�g�m�G��I����V��_�D��d�d�e�e�u�}�W���[����V��^�D��d�e�d�d�f�l�F��I����FǻN��E��e�e�e�e�g�m�G��I����W��_�E��y�_�u�u�g�m�G��I����V��^�D��d�d�e�e�g�l�[�ԜY���V��^�E��d�e�e�e�f�l�F��I����W�d��U���e�e�e�e�g�l�G��H����W��_�D��e�w�u�u�w��G��I����W��_�E��d�d�d�d�f�l�F���Y���D��^�E��e�d�d�e�g�m�F��H����V��L����u�e�e�e�g�m�F��I����W��_�D��d�e�d�y�]�}�W��I����V��^�E��d�d�d�d�f�m�F��H���F�^�E��e�e�e�d�f�l�G��H����V��_�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�d�u�}�W���[����V��^�D��d�e�e�d�f�l�F��H����FǻN��E��e�e�e�d�f�l�F��I����W��_�D��y�_�u�u�g�m�G��I����V��_�D��d�d�d�e�g�l�[�ԜY���V��^�E��d�d�e�e�f�l�F��H����W�d��U���e�e�e�e�g�l�G��H����W��_�E��e�w�u�u�w��G��I����W��_�D��d�d�d�d�g�l�G���Y���D��^�E��d�e�e�d�g�m�F��H����W��L����u�e�e�e�g�m�F��H����W��_�D��e�d�d�y�]�}�W��I����V��^�D��d�d�d�d�f�l�G��H���F�^�E��e�e�d�e�f�l�G��H����W��^�W���u�u�w�e�g�m�G��H����W��_�D��d�e�e�e�u�}�W���[����V��^�D��e�e�d�d�f�l�F��I����FǻN��E��e�e�e�d�f�m�G��I����W��^�E��y�_�u�u�g�m�G��I����W��_�D��d�d�d�d�f�m�[�ԜY���V��^�E��d�d�d�e�f�l�F��H����V�d��U���e�e�e�e�f�m�G��H����W��_�D��e�w�u�u�w��G��I����V��_�E��d�d�d�d�f�m�G���Y���D��^�E��e�e�d�e�g�l�F��H����V��L����u�e�e�e�g�m�G��H����V��_�D��e�e�d�y�]�}�W��I����V��^�D��d�d�d�d�f�l�G��H���F�^�E��e�d�e�d�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�d�e�e�u�}�W���[����V��_�E��d�d�e�d�f�l�F��I����FǻN��E��e�e�e�e�g�m�G��I����W��_�D��y�_�u�u�g�m�G��I����V��^�D��d�d�d�d�g�m�[�ԜY���V��^�D��d�d�e�d�f�l�F��H����V�d��U���e�e�e�e�f�m�F��H����W��_�D��e�w�u�u�w��G��I����V��_�E��d�d�d�d�f�l�F���Y���D��^�E��e�e�e�d�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�d�e�y�]�}�W��I����V��^�D��e�e�e�e�g�m�G��I���F�^�E��e�d�e�d�f�l�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�d�u�}�W���[����V��_�E��d�e�d�e�g�m�G��H����FǻN��E��e�e�e�e�g�m�G��H����V��^�D��y�_�u�u�g�m�G��I����W��^�E��e�e�e�d�g�l�[�ԜY���V��^�D��e�d�e�e�g�m�G��I����W�d��U���e�e�e�e�f�m�G��H����V��^�E��e�w�u�u�w��G��I����V��_�D��e�e�e�e�g�m�F���Y���D��^�E��e�e�e�d�f�m�G��I����W��L����u�e�e�e�g�m�G��I����V��^�E��d�e�e�y�]�}�W��I����V��_�D��d�e�e�e�g�m�F��I���F�^�E��e�e�d�d�g�l�G��I����V��_�W���u�u�w�e�g�m�G��H����W��^�E��e�e�d�d�u�}�W���[����V��^�D��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�d�f�l�G��H����V��_�E��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�f�m�[�ԜY���V��^�E��e�e�d�e�g�m�G��I����W�d��U���e�e�e�e�g�l�F��I����V��^�D��d�w�u�u�w��G��I����W��^�D��e�e�e�e�f�l�G���Y���D��^�E��d�e�e�e�f�m�G��I����W��L����u�e�e�e�g�m�F��H����V��^�E��e�e�e�y�]�}�W��I����V��^�E��d�e�e�e�g�m�G��I���F�^�E��e�e�d�e�f�m�F��I����V��_�W���u�u�w�e�g�m�G��I����V��^�E��e�d�d�d�u�}�W���[����V��^�D��e�d�e�e�g�m�G��H����FǻN��E��e�e�e�d�f�m�F��I����V��_�D��y�_�u�u�g�m�G��I����W��_�E��e�e�e�d�g�m�[�ԜY���V��^�E��e�d�e�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��I����V��^�D��d�w�u�u�w��G��I����V��^�E��e�e�e�e�f�m�F���Y���D��^�E��d�e�e�d�f�l�G��I����V��L����u�e�e�e�g�m�F��H����W��^�E��d�e�d�y�]�}�W��I����V��^�D��e�e�e�e�g�m�F��I���F�^�E��e�e�e�e�g�m�G��I����V��_�W���u�u�w�e�g�m�G��H����W��^�E��e�d�e�e�u�}�W���[����V��^�D��d�e�d�e�g�m�G��I����FǻN��E��e�e�e�e�f�l�G��I����V��_�D��y�_�u�u�g�m�G��I����V��^�E��e�e�e�d�f�l�[�ԜY���V��^�E��d�d�d�e�g�m�G��I����W�d��U���e�e�e�e�g�l�F��H����V��^�D��e�w�u�u�w��G��I����W��^�E��e�e�e�e�f�m�G���Y���D��^�E��e�e�d�d�f�m�G��I����V��L����u�e�e�e�g�m�G��I����W��^�E��d�d�d�y�]�}�W��I����V��_�D��e�e�e�e�g�m�F��I���F�^�E��e�e�e�d�g�m�G��I����V��_�W���u�u�w�e�g�m�G��I����W��^�E��e�d�e�e�u�}�W���[����V��^�D��d�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�f�m�G��H����V��_�E��y�_�u�u�g�m�G��I����W��_�E��e�e�e�d�g�l�[�ԜY���V��^�E��d�e�e�d�g�m�G��I����V�d��U���e�e�e�e�g�m�F��I����V��^�D��e�w�u�u�w��G��I����V��_�E��e�e�e�e�f�m�G���Y���D��^�E��e�e�e�d�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��d�e�e�y�]�}�W��H����W��_�E��e�e�e�e�g�m�G��H���F�_�D��d�d�d�d�f�m�F��I����V��_�W���u�u�w�d�f�l�F��H����V��^�E��e�d�d�e�u�}�W���[����W��_�D��e�e�e�e�g�m�G��H����FǻN��D��d�d�d�d�f�m�F��I����V��_�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�e�g�l�[�ԜY���W��_�D��d�e�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�D��e�w�u�u�w��F��H����W��_�E��e�e�e�e�f�l�G���Y���D��_�D��d�e�d�d�g�l�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�d�e�y�]�}�W��H����W��^�E��e�e�e�e�g�m�G��I���F�_�D��d�d�e�d�f�m�F��I����V��^�W���u�u�w�d�f�l�F��I����V��^�E��e�d�e�d�u�}�W���[����W��_�D��e�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��H����V��_�E��y�_�u�u�f�l�F��H����W��_�E��e�e�e�d�f�l�[�ԜY���W��_�D��e�e�e�d�g�m�G��I����V�d��U���d�d�d�d�f�m�G��H����V��^�E��e�w�u�u�w��F��H����V��^�D��e�e�e�e�g�l�F���Y���D��_�D��d�e�d�d�f�l�G��I����W��L����u�d�d�d�f�l�F��H����V��^�E��d�e�d�y�]�}�W��H����W��^�E��e�e�e�e�g�m�F��H���F�_�D��d�d�e�d�f�l�F��I����V��_�W���u�u�w�d�f�l�F��I����W��^�E��e�e�e�e�u�}�W���[����W��_�E��e�d�e�e�g�m�G��I����FǻN��D��d�d�d�d�g�l�F��I����V��^�E��y�_�u�u�f�l�F��H����W��^�E��e�e�e�d�g�l�[�ԜY���W��_�D��e�e�e�d�g�m�G��I����V�d��U���d�d�d�d�f�m�G��I����V��^�E��d�w�u�u�w��F��H����V��_�D��e�e�e�e�g�l�G���Y���D��_�D��d�e�e�e�g�l�G��I����W��L����u�d�d�d�f�l�F��I����V��^�E��e�e�d�y�]�}�W��H����W��^�E��d�e�e�e�g�m�G��I���F�_�D��d�d�e�e�g�l�F��I����V��^�W���u�u�w�d�f�l�F��I����V��^�E��e�e�e�d�u�}�W���[����W��_�E��e�e�d�e�g�m�G��I����FǻN��D��d�d�d�e�f�l�F��I����V��^�D��y�_�u�u�f�l�F��H����W��^�E��e�e�e�e�f�m�[�ԜY���W��_�D��d�d�e�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�G���Y���D��_�D��e�d�d�d�f�l�F��H����W��L����u�d�d�d�f�l�G��H����W��_�D��d�d�e�y�]�}�W��H����W��_�D��d�d�d�d�f�l�F��H���F�_�D��d�d�d�d�f�l�F��H����W��_�W���u�u�w�d�f�l�F��I����V��_�D��d�d�d�d�u�}�W���[����W��_�E��e�e�e�d�f�l�F��H����FǻN��D��d�d�d�d�g�m�F��H����W��_�E��y�_�u�u�f�l�F��H����V��^�D��d�d�d�d�g�m�[�ԜY���W��_�D��e�d�e�d�f�l�F��H����W�d��U���d�d�d�d�f�m�G��H����W��_�D��d�w�u�u�w��F��H����V��_�D��d�d�d�d�f�m�G���Y���D��_�D��d�e�d�e�g�m�F��H����V��L����u�d�d�d�f�l�F��H����V��_�D��d�d�e�y�]�}�W��H����W��^�E��e�d�d�d�f�l�F��H���F�_�D��d�d�e�e�f�l�F��H����W��^�W���u�u�w�d�f�l�F��I����W��_�D��d�d�e�e�u�}�W���[����W��_�E��e�e�e�d�f�l�F��I����FǻN��D��d�d�d�d�g�m�F��I����W��_�E��y�_�u�u�f�l�F��H����V��^�D��d�d�d�e�f�l�[�ԜY���W��_�D��d�d�d�d�f�l�F��H����W�d��U���d�d�d�d�f�m�F��H����W��_�D��d�w�u�u�w��F��H����V��^�D��d�d�d�d�f�l�G���Y���D��_�D��d�e�d�d�g�m�F��H����W��L����u�d�d�d�f�l�F��I����V��_�D��e�d�e�y�]�}�W��H����W��_�E��d�d�d�d�f�l�G��I���F�_�D��d�d�e�e�f�l�F��H����W��^�W���u�u�w�d�f�l�F��I����V��_�D��d�d�d�d�u�}�W���[����W��_�D��d�e�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�l�G��I����W��_�E��y�_�u�u�f�l�F��H����V��_�D��d�d�d�e�g�m�[�ԜY���W��_�D��d�e�d�d�f�l�F��H����V�d��U���d�d�d�d�f�m�F��I����W��_�D��e�w�u�u�w��F��H����V��^�E��d�d�d�d�f�l�G���Y���D��_�D��d�d�d�d�f�l�F��H����W��L����u�d�d�d�f�l�F��H����V��_�D��e�e�d�y�]�}�W��H����W��^�E��d�d�d�d�f�l�G��H���F�_�D��d�d�d�e�f�m�G��H����W��^�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�e�u�}�W���[����W��_�E��d�d�e�d�f�l�F��H����FǻN��D��d�d�d�d�g�l�G��I����W��_�E��y�_�u�u�f�l�F��H����V��_�D��d�d�d�e�g�m�[�ԜY���W��_�D��d�e�d�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��I����W��_�D��e�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�G���Y���D��_�D��d�e�d�e�g�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��e�e�d�y�]�}�W��H����W��_�E��e�d�d�d�f�l�G��H���F�_�D��d�d�d�e�f�m�F��H����W��^�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�e�u�}�W���[����W��_�D��d�d�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�l�G��H����W��_�E��y�_�u�u�f�l�F��H����V��^�D��d�d�d�e�g�m�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��H����W��_�D��d�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�d�d�f�l�F��H����W��L����u�d�d�d�f�l�F��H����V��_�D��e�e�d�y�]�}�W��I����V��^�E��e�d�d�d�f�l�G��I���F�^�E��e�e�e�e�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�d�d�e�u�}�W���[����V��^�E��d�e�e�d�f�l�F��H����FǻN��E��e�e�e�e�g�l�G��H����W��_�D��y�_�u�u�g�m�G��I����W��_�D��d�d�d�e�f�m�[�ԜY���V��^�E��e�d�e�e�f�l�F��H����V�d��U���e�e�e�e�g�m�F��I����W��_�D��d�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�F���Y���D��^�E��e�e�e�e�g�l�F��H����V��L����u�e�e�e�g�m�G��I����W��_�D��d�e�e�y�]�}�W��I����V��^�E��d�d�d�d�f�l�F��H���F�^�E��e�e�e�d�g�m�G��H����W��^�W���u�u�w�e�g�m�G��I����V��_�D��d�d�e�d�u�}�W���[����V��^�E��e�d�d�d�f�l�F��I����FǻN��E��e�e�e�e�g�l�F��H����W��_�E��y�_�u�u�g�m�G��I����V��_�D��d�d�d�d�g�l�[�ԜY���V��^�E��e�e�e�e�f�l�F��H����V�d��U���e�e�e�e�g�m�G��H����W��_�D��e�w�u�u�w��G��I����V��_�E��d�d�d�d�f�m�G���Y���D��^�E��e�d�e�d�f�l�F��H����V��L����u�e�e�e�g�m�G��I����W��_�D��d�d�e�y�]�}�W��I����V��_�E��e�d�d�d�f�l�F��H���F�^�E��e�e�e�e�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�e�u�}�W���[����V��^�D��e�e�e�d�f�l�F��H����FǻN��E��e�e�e�e�f�l�G��H����W��_�E��y�_�u�u�g�m�G��I����W��^�D��d�d�d�d�g�l�[�ԜY���V��^�E��e�d�e�d�f�l�F��H����V�d��U���e�e�e�e�g�m�G��H����W��_�D��d�w�u�u�w��G��I����V��^�E��d�d�d�d�f�l�F���Y���D��^�E��e�d�e�e�f�l�F��H����W��L����u�e�e�e�g�m�G��I����W��_�D��d�d�e�y�]�}�W��I����V��_�E��e�d�d�d�f�l�F��I���F�^�E��e�e�e�d�g�m�G��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�d�d�e�u�}�W���[����V��^�D��d�d�d�d�f�l�F��H����FǻN��E��e�e�e�e�f�m�F��I����W��_�D��y�_�u�u�g�m�G��I����V��_�D��d�d�d�d�f�l�[�ԜY���V��^�E��d�e�d�e�f�l�F��H����W�d��U���e�e�e�e�g�m�F��H����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�d�e�d�f�l�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�d�y�]�}�W��I����V��_�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�d�g�m�F��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�d�u�}�W���[����V��^�D��e�d�d�e�g�m�G��I����FǻN��E��e�e�e�e�f�m�G��H����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�f�m�[�ԜY���V��^�E��d�e�e�d�g�m�G��I����V�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��_�E��e�e�e�e�g�m�G���Y���D��^�E��e�d�d�d�f�m�G��I����V��L����u�e�e�e�g�m�G��H����W��^�E��e�d�d�y�]�}�W��I����V��_�D��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�f�m�F��I����V��_�W���u�u�w�e�g�m�G��I����W��^�E��e�e�e�d�u�}�W���[����V��^�D��d�d�d�e�g�m�G��I����FǻN��E��e�e�e�e�f�l�F��I����V��^�D��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�f�l�[�ԜY���V��^�E��e�e�e�d�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�E��d�w�u�u�w��G��I����V��_�E��e�e�e�e�g�m�F���Y���D��^�E��e�d�e�e�f�m�G��I����W��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��_�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�e�u�}�W���[����V��^�D��e�e�d�e�g�m�G��H����FǻN��E��e�e�e�e�g�l�F��H����V��^�E��y�_�u�u�g�m�G��I����W��^�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�d�d�e�g�m�G��I����W�d��U���e�e�e�e�g�m�F��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�l�G���Y���D��^�E��e�e�d�e�f�l�G��I����W��L����u�e�e�e�g�m�G��H����V��^�E��e�e�d�y�]�}�W��I����V��^�D��e�e�e�e�g�m�G��H���F�^�E��e�e�e�d�f�m�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��H����FǻN��E��e�e�e�e�g�m�F��H����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�l�[�ԜY���V��^�E��d�e�d�e�g�m�G��I����W�d��U���e�e�e�e�g�m�G��H����V��^�E��e�w�u�u�w��G��I����V��_�D��e�e�e�e�g�l�G���Y���D��^�E��e�e�d�e�f�l�G��I����W��L����u�e�e�e�g�m�G��H����W��^�E��e�e�d�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����W��^�E��e�e�d�e�u�}�W���[����V��^�E��e�d�e�e�g�m�G��H����FǻN��E��e�e�e�e�g�m�F��H����V��^�E��y�_�u�u�g�m�G��I����V��_�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�d�d�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�D��e�e�e�e�g�l�G���Y���D��^�E��e�e�e�d�f�l�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�d�d�y�]�}�W��I����V��^�E��d�e�e�e�g�m�G��H���F�^�E��e�e�e�e�g�m�G��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�d�u�}�W���[����W��_�D��d�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�l�G��I����V��^�D��y�_�u�u�f�l�F��H����W��_�E��e�e�e�e�f�m�[�ԜY���W��_�D��d�d�e�e�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��d�w�u�u�w��F��H����W��^�D��e�e�e�e�g�m�F���Y���D��_�D��d�d�d�e�f�l�G��I����V��L����u�d�d�d�f�l�F��H����V��^�E��e�d�d�y�]�}�W��H����W��_�E��e�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�m�G��I����V��_�W���u�u�w�d�f�l�F��H����W��^�E��e�e�e�e�u�}�W���[����W��_�D��d�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��H����V��^�D��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�f�m�[�ԜY���W��_�D��d�d�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��_�D��e�e�e�e�g�m�F���Y���D��_�D��d�d�e�e�g�l�G��I����V��L����u�d�d�d�f�l�F��I����V��^�E��e�e�d�y�]�}�W��H����W��_�E��d�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�d�u�}�W���[����W��_�D��d�e�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�F��H����V��^�E��y�_�u�u�f�l�F��H����V��^�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�d�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��H����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�e�g�m�G��I����V��L����u�d�d�d�f�l�F��I����W��^�E��e�e�d�y�]�}�W��H����W��_�E��e�e�e�e�g�m�G��H���F�_�D��d�d�d�d�g�l�G��I����V��^�W���u�u�w�d�f�l�F��H����V��^�E��e�e�e�e�u�}�W���[����W��_�D��e�d�d�e�g�m�G��I����FǻN��D��d�d�d�d�f�m�G��H����V��^�E��y�_�u�u�f�l�F��H����V��_�E��e�e�e�e�g�m�[�ԜY���W��_�D��d�e�e�d�g�m�G��I����V�d��U���d�d�d�d�f�l�F��I����V��^�E��e�w�u�u�w��F��H����W��^�E��e�e�e�e�g�m�G���Y���D��_�D��d�d�e�e�g�m�F��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�d�y�]�}�W��H����W��_�E��d�d�d�d�f�l�F��H���F�_�D��d�d�d�d�g�l�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�D��e�d�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��I����W��_�D��y�_�u�u�f�l�F��H����V��^�D��d�d�d�d�f�l�[�ԜY���W��_�D��d�e�e�e�f�l�F��H����V�d��U���d�d�d�d�f�l�F��I����W��_�D��d�w�u�u�w��F��H����W��^�D��d�d�d�d�f�l�F���Y���D��_�D��d�d�e�d�f�m�F��H����W��L����u�d�d�d�f�l�F��I����V��_�D��d�d�e�y�]�}�W��H����W��_�E��d�d�d�d�f�l�F��I���F�_�D��d�d�d�d�g�l�G��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�D��e�e�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�G��H����W��_�D��y�_�u�u�f�l�F��H����V��_�D��d�d�d�d�f�m�[�ԜY���W��_�D��d�d�e�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��H����W��_�D��d�w�u�u�w��F��H����W��_�D��d�d�d�d�f�l�F���Y���D��_�D��d�d�e�e�f�l�F��H����W��L����u�d�d�d�f�l�F��I����W��_�D��d�d�e�y�]�}�W��H����W��_�D��d�d�d�d�f�l�F��I���F�_�D��d�d�d�d�f�m�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�e�u�}�W���[����W��_�D��d�e�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�m�F��I����W��_�D��y�_�u�u�f�l�F��H����W��^�D��d�d�d�d�f�l�[�ԜY���W��_�D��d�e�e�d�f�l�F��H����W�d��U���d�d�d�d�f�l�F��I����W��_�D��e�w�u�u�w��F��H����W��^�E��d�d�d�d�f�l�G���Y���D��_�D��d�d�d�e�g�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�d�y�]�}�W��H����W��_�E��d�d�d�d�f�l�F��I���F�_�D��d�d�d�d�g�m�F��H����W��_�W���u�u�w�d�f�l�F��H����V��_�D��d�d�d�d�u�}�W���[����W��_�D��d�d�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�l�F��H����W��_�D��y�_�u�u�f�l�F��H����W��^�D��d�d�d�d�f�m�[�ԜY���W��_�D��d�e�d�d�f�l�F��H����V�d��U���d�d�d�d�f�l�F��I����W��_�D��d�w�u�u�w��F��H����W��_�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�d�e�f�l�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�e�y�]�}�W��H����W��_�D��e�d�d�d�f�l�F��I���F�_�D��d�d�d�d�f�l�F��H����W��_�W���u�u�w�d�f�l�F��H����W��_�D��d�d�d�d�u�}�W���[����W��_�D��e�d�d�d�f�l�F��H����FǻN��D��d�d�d�d�f�l�F��H����W��_�D��y�_�u�u�f�l�F��H����W��^�D��d�d�d�d�f�m�[�ԜY���W��_�D��d�d�e�e�f�l�F��H����V�d��U���d�d�d�d�f�l�F��I����W��_�D��d�w�u�u�w��F��H����W��_�E��d�d�d�d�f�l�F���Y���D��_�D��d�d�d�d�g�m�F��H����W��L����u�d�d�d�f�l�F��H����W��_�D��d�d�e�y�]�}�W��H����W��_�D��e�d�d�d�f�l�F��I���F�_�D��d�d�d�d�f�l�F��H����W��_�W���u�u�w�e�g�m�G��I����V��_�D��d�d�d�d�u�}�W���[����V��^�E��e�e�d�d�f�l�F��H����FǻN��E��e�e�e�e�g�m�G��H����W��_�D��y�_�u�u�g�m�G��I����V��_�D��d�d�d�d�f�l�[�ԜY���V��^�E��e�e�e�e�f�l�F��H����W�d��U���e�e�e�e�g�m�G��I����W��_�D��d�w�u�u�w��G��I����V��^�D��d�d�d�d�f�l�F���Y���D��^�E��e�e�e�e�g�m�F��H����W��L����u�e�e�e�g�m�G��I����W��_�D��d�d�d�y�]�}�W��I����V��^�E��d�d�d�d�f�l�F��H���F�^�E��e�e�e�e�g�l�F��H����W��_�W���u�u�w�e�g�m�G��I����W��_�D��d�d�d�d�u�}�W���[����V��^�E��e�d�d�d�f�l�F��H����FǻN��E��e�e�e�e�g�m�G��H����W��_�D��y�_�u�u�g�m�G��I����V��_�D��d�d�d�d�f�l�[�ԜY���V��^�E��e�e�d�d�f�l�F��H����W�d��U���e�e�e�e�g�m�G��H����W��_�D��d�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�d�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��d�e�d�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�F��H����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�d�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�d�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��d�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��L����u�e�e�e�g�m�G��I����V��^�E��e�e�e�y�]�}�W��I����V��^�E��e�e�e�e�g�m�G��I���F�^�E��e�e�e�e�g�m�G��I����V��^�W���u�u�w�e�g�m�G��I����V��^�E��e�e�e�e�u�}�W���[����V��^�E��e�e�e�e�g�m�G��I����FǻN��E��e�e�e�e�g�m�G��I����V��^�E��y�_�u�u�g�m�G��I����V��^�E��e�e�e�e�g�m�[�ԜY���V��^�E��e�e�e�e�g�m�G��I����V�d��U���e�e�e�e�g�m�G��I����V��^�E��e�w�u�u�w��G��I����V��^�E��e�e�e�e�g�m�G���Y���D��^�E��e�e�e�e�g�m�G��I����V��LךU���x�z��&��8������ƹF�N�����4�>�2�u��:����0����C%��Q�����&�_�_