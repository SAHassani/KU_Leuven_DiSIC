-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B/��B�����;�g�6�#�3�p�W�������w��u�����u�'�2�;�;������Ɯ�z��Z������!�o�d�w�<����Y����9K��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�w�>�W��Jӥ��J��_�����;�9��&�%�0����:����A��X חXʔ�9��2�!�w�8�������}��X ��U���!� �0�!�w�3����ӯ��\��C�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z��Y����\��=C�Uʁ�<�u�:�%�9�3�W�������G��^ ��ʦ�8�9�;�{�w�2�W���Ӕ��\��RN�����4�<�;�x�w�}��������F��R�����#�'�<�;�w�;����Y����\��CN��ʾ�#�'�9�6�]�p�Wϻ�����F��SN�Uʚ�=�'�#�9�2�}�����ƿ�C��C�����=�&�!�8�y�p�}��YӲ��@F��Z�����!�>�&�<�w�����Y����@"��V8�����y�4�1�%�8�(��ԑT����@"��V=�����y�&��!��1����	�����������<�{�u�&�6�<�����ƭ�G��[חX���6�8�&�<�w�*�W�������@"��V(�����8�9�1�4�3�.�3���*����W5��G��[���=�_�x�u�u�4�����Ƹ�VF��X��U���2�0�0�!�w�3�W���Yѕ��\�������,�1�7�u�9�W�Z�������R
��V�����u�,�9�{�w�5�����ƹ�V��V��U�����7��#�/��������[ǶN��8����4�;�!�2�9�����Ʃ�R��DN�����9�u�9�2�2�q����Ӊ��D��_N��ʳ�9�0�_�x�w�4�W���s��ƴF�D�� ���0�u�&� �2�}����Y����A��RN��ʦ��1��4�9�}�Ϫ�Ӓ����Z���߇x�u� �0�w�3��������_�CחX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�W�����ƥ�V��N��ʼ�0�{�!�
�8�4�(��M݇��l�B�����{� �0�<��)�Y���B���Q��NN����u� �0�"�%�s����W����9F��D������2�<�!�;�)����	݇��l��Y��ʐ��%�!�4�'�4�ݱ�Y����V��^��Uʾ�4�4�<�!�w�}�W���Y����]F��C��ʧ�;�0�d�u�8�l�W��H��ƹ��TN��U���u�u�u�u�w�}�Ϸ�������P��U���d�u�o�u�w�f����Q����R��R-��;���u�u�u�u�w�3��������lǻ������6�u�u�w�}�W���ӥ��]��T1�����&�4�4�4�>��W���Y�����D�����6�_�u��#��W���Y���F�N��U����!�
�}��>�FϺ�����O��N��1����'�!�4�'�8�W������C��C��]���6�d�1�"�#�}�^��Yۉ��V��	F�����h�r�r�|�]�}��������]��Z����:�!��6�6�<�ǵ�	����W	��C��\��u�:�=�'�j�u����
���O�=N�����4�4�<��:�1����Y����@��[�����6�:�}��4�l��������\������k�e�|�_�w�.�������F�N��Oʺ�!�&�1�9�0�>�M���I���9��+������8�9�;�e�>�}�������V��E��!���3���%�#�<��������ZǑN����>�&�2�!�%�W�W�������@��Y
װUʶ�;�!�;�u��8�������\��Y�����4�2�u�u�8�n�M���B���K��_��U���4�&�4�0�6�.����ӂ��RF��G��ʰ�&�'�u�;�.�)�ϫ��Ʈ�G��EךU���<�6� �0�w�3����[����F��C�� ���u��r�u�>�8�ϭ�������YN��ʻ�'�4�_�u�z���������J��=N�����u��4�9�6�<����&�ƥ���V�����x�u�:�;�8�m�W���
����\��h�����>�4�4�<�#�p�W������]ǻ�����&��!��2�}�W���Y�Ɵ�R
��V�����
�u�h�}�#�8��������@[�I��N�ߊu�<�;�9�$���������V�N�����2�6�#�6�8�u�$���Hӂ��]��G��H���!�0�&�k�g�t�}���������V������,�u�o�$�9��������G	��\=��X���:�;�:�e�w�`�_������V�dךU���;�9�&��#�����Y���	F��V�����'�4�
�u�j�u����
����G��DS�E���n�u�&�2�6�}��������]�N��U���9��!��%�$���Yۉ��V��	F�����h�r�r�|�]�}�����ƿ�d��V�����u�u�u�!��2����D����lǻ�����&�� �!�2�����Y�Ǝ�\
��Y8�����>�%�x�u�8�3���Y���\��E�����0�n�_�u�z�����Ӓ�� ����U���4�<�y�!�w�+��������V�������"�!�u�=�w�)��ԜY����z4��_�� ���u�=�&�&�:�}����Q����[��fN�����{�u�4�!�>�(�ϵ�����@��Y	�Uʴ�!�<� �0�<�8�W���
����R>��EN��U���u�o�&�2�6�}�������9F��C�����u�0�%�:�w�.��������U��N��U���;�9�<�u�#�(�U�ԜY����Z��RN�����3�&�� �#�8�2������	F��P ��U���w�'�0�n�w�<��������V��X�����=�<��9�w�}�W��
����_F��L�� ���_�u�!�'�5�)�W���	Ӊ��@��C�����u�u�u�u�w�4��������A��d�����<� �0�>�2�}�ϭ�=����V��SN��U���o�&�2�4�w�.�U�����ƓF�:��U���<�&�:�u�?�}��������@F��E�����8�;�1�0�'�/����������[�����u�x�u�=�8�:�W�������G��Y	�����!�_�u�!�%�?��������]	��N�����n�u�4�!�>�(�ϳ�����\��X�����=�<��9�m�.����Y���D��N����� �0�8�-�1�3����ӕ��R��^��U��&�2�4�u�$��U�ԜY����Z��RN�����;� �u�3�$���������	F��P ��U���w�w�_�_�]�8��ԶY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x��%�!��0����s���F�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߊu�x��0�2�4�W�������V��[�����u�3�&��#��[ϭ�=����R
��~ �����4�;�e�{�}�Z����ƿ�r��t����u�&�!�0�w�/�W����Ƽ�@����U���!�<�u�:�'�3�������K��Y�����0�&�7�<�#�/�Wϭ�=����]F��X��U���9�;�1� �w�4�ϭ�8����[��^�E�ߊu�x�&��#�����ӕ��F
��G�����<�u�,�:�2�.����UӇ����R-�����|�&�:�9�]�}�ZϮ�������U�����0�u�4�%�2�}�#���Y����Z��V��ʡ�4�u�=�"�w�3�W��Y����A�\��ʡ�0��9�;�w�4����MӢ����EN�����}�2�b�{�3�}�Ϯ�����VO�N�U���u�=�u�9�0�0����
ӕ��T��R
�� ���:��&�!�6�}��������R��SN�����'�4�_�u�z�)�W�������G��Y	�U���_�u�x�u�z�}��������P
��\S�U���u�u�u�u�w�}�W���Y����l9�N��*���u�u�
�u�w�}�(���Y�Ɠ�lF�N��*���u�
�
�u�z�}���������N��	���)�
�)�u�+���������F��h1��U���
�
�u�u���W���&���KǻC����1��4�;�g�}�WϢ�Y����^��U���u�u�u�u�w�}�W���Y���OF�N��	���d�u�_�u�z�}�W���Y���F�1��*���
�
�
�
���(���&����l9��h1��*���
�u�
�
���(���&���F��s��<���'�!�u�
���(�������l9��1��*���
�
�
�u�w��(���&����lF��h1��*�ߊu�x�u�u�w�}�W���Y����l9��h1��*���
�
�
�u�w�}�W���Y���9��h1��*���
�
�
�
���W��Y����G��[�����u�u�u�u�w�}�W���YӚ��l9��h1��*���
�_�u�x�w�}�W���Y���F�N��U���u�
�
�
��}�W���Yӹ��l9��N��U���u�
�
�
�]�}�Zϭ�.����Z�N��U���
�
�
�
�w�}�W���&����l9��N��Uʩ�
�
�
�)�w�}�WϢ�&����9F�d��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}��������^��d�����0�&��8�;�����s�Ʈ�T��N�����<�<�2�0�0�u��������KO��_�����u�u�:�u�w�3�GϪ�Y����W��X��U���u�u�x�u�%�<�Ͽ�?�ƺ�A��YN��U���&�:�0�6�4�8���� Ӏ����^ ��U���u�u�&��"�)��������zO�
N��6���!�0�}�|�u�m�L�ԜY���F�:������u�'�;�1�/����Y������X��ʡ�u�=�u�-�3�0���Y����VF��Rd��U���u�x�u�0�'�}�Ϫ��Ƹ���B�����u�:�r�u�2�}����ӑ��[F��G�����u�;�u�u�w�}�Z�������u/�������!�0��{�w�}�W����ƿ�p	��C8��0���9�}�|�!�2�W�W���Y���@��C�����|�>�4�4�>�)�Z�������V�S��1����}�|�>�6�<����T�ƨ�D��^����u�u�u�u�$�<��������AN��R�����4�4�<��l�}�W���YӃ����=d��U���u�x�u�0�3�)�W����Ƹ�VF��C�����8�9��<�>����Y����]��Y����� �!�u�u�w�}�Z����ƨ�G��[�����4�{�u�=�$�4�W���Ӏ����L�����u� �%�!�]�}�W���Y����@"��V8�����0�}�|�r�p�<�ϭ�:����e��F��D�u�=�;�u�w�}�W���
����R ��D��\��u�&�4�4�1�/�>��Y���F��Y
���ߠu�u�u�u�>�}��������v��[_��\ʡ�0�_�u�u�w�}�W�������P	��'��I���&�4�4�<�$�u�^�ԜY���F��SN��N�ߊu�u�u�;�w�2��ԶY�����V������,�i�u�$�<��������A]ǑN��U���u�0�=�<��}���� ����Q��E�����4�<�_�u�w�}�ϭ�:����e��G��:���6�:�>�d�#�8�}���Y���@��t�����u�h�r�r�w�1�ϭ�.����Z��[N�U��n�u�u�u�2�9���s���V��^�X���<�<�2�0�0�W�W���Y����V��g��!����8�<�n�]�}�Z�������@��[��U���u�:�0�"�#�}����Y������RN�����=�u�<�=�w�4����ӄ��@��=N��Xʢ�u�<�;�!�u�8�����Ʃ�G��q(��[���:�0�0�u�?�}����?����AF��G��U���_�u�x� �>�:����*����G�������=�6�u�:�$�z�W���Ӎ��G��S��Uʆ�u�0�<�0�#�W�W��������C@��!���0�0�!�4�g�.� ���Y����C��^��U���u�!�6�8�>�8����W���a��M�����'�!�u�'�4�.�_�������A��=N�����_�u�u�&�6�<����*����V�
N�����&�k�:�=�%�`�P���P���F��EN�����u�:�>�%�z�}����Y�����V������8�9�1��u�3���.����W��X����u�h�&��#�����0��ƹF��Y
�����_�u�;�u�%�>��������w��q���ߠu��&�/��)�$�������A	��D�����4�0�:�1�]�}����s���@��C������8�9�1�k�}�������\��E��R��|�_�u�u�8�}�W���IӒ��X5��_�����u�u�u�&��)�$�������C
��'�����4�<�!�x�w�2����I�����V�����1��n�u�w�8�ϲ���ƹ�������u�0�<�0�6�<������ƓF��`�����i�u�&�0�?�4�;���s�ƿ�w��a�����%�0�u�h�$���������J]ǑN�U���u�3��%�#��������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�0�1���W