-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B%��Q"�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������4ǶN����g�u�4� �%�}�G��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�6�u�g�l�4�������(��^��ʜ�&�'�8�;�$���������9K�v��'���!�u�0�0�!�9�Z�������R
��Y�� ���!�u�;�0�9�1�>�������\ǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x�z�}����
����[��T�����!�!�>�&�>�}��������P��CN�����<�;�9�y�6�9��������K������ �9�&�2�6�.��������\ ��_��4���u��0�6�2�;�����Ƣ�V��XN��U���u�u�:�1�3�4�W���	����_F��S��U���u�=�u�:�2�}�ϛ�*����V ��C�����8�'�u�;�8�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�Cװ���'�'�u�0�2�W�W���Y������h�����d�a�4�9�]�}��������F��^�����9�n�_�;�>�$�2�������W��^�����0�<�}�u�<�+�������F��^ �����0�u�h�f�]�}�4���.����F�T��ʼ�!�2�'�o�w�e�}���7����P�N��U���;�<�!�2�%�g�W��P���A�N������>�u�u�w�}�ϭ�����Z��N������>�-�u�w�}�ϭ�����Z��=N��6����4�u�u�w�g��������T��=N��6����u�u�u�w�g��������T��=N��6����;�u�u�w�g��������T��A������0��1�?�l��������lǻ�����1�'�u�u�m�2�ϭ�����Z��R����1�"�!�u�~�W�W�������r��NN��U���u�!�
�:�>�����ۍ��^+��DC����!�u�|�_�w�.�������F���U���
�:�<�
�2�)�ǵ�����W��N�����u�|�_�u�$�2����:����\��B�����:�<�
�0�#�/����4����F��@ ��U���|�_�;�u�&�2��������9l��T�����'�u��u�1��4���5����AF��=d��X���<�6�u�=�%�}��������X5�������0��0�u�8�9����Ӓ�� ��[N��U���!�'�u�u�z�}��������@F���� ���!�0�u�:�p�}����������R��ʴ�1�6� �0�#�0����
����9F��^	��ʦ�:�3�:�1�2�}�W���Cӕ��l
��^��H��r�_�u�<�9�1��������TF�N��U���!�
�:�<�w�`�P���s�ƿ�T�������;�0�u�u�w�}�W���&����P9��T��]���0��1�=�f�9� ���Y���F��C����e�|�_�u�>�3�ϭ�����F��EN��U���u�;�<�;�3�l��������\������k�e�|�_�w�4����
����Z ��N��U���u�u�!�
�8�4�(�������}��V��Dʱ�"�!�u�|�m�}�������A�=N�����9�&��0��9�;���Y�����h�����0�!�'�d�3�*����P���	��R��K��|�_�u�<�9�1��������p	��D"��U���!�
�:�<��8��������R��N�����u�|�o�u�8�5���^���9F��^	��ʦ��0��!��1�W���Cӕ��l
��^�����'�>�:�3�>�)�Z�������V�S�����'�h�r�r�l�}�����ƿ�p	��`�����6�u�o�&�3�1��������AN��B�����u�:�;�:�g�}�J�������X�G�Uʦ�2�4�u�&�8�;����Y���F��D�����6�o�u�e�l�}�����ƿ�p	��`�����u�u�o�&�3�1����C���]ǑN����� �0�>�0�w�}�������R��^��ʾ�0�u�3�&�8�;�������F��D�����&�w�'�0�l�}����������GN��U���0���2�w�}�W��
����_F��L�� ���_�u�!�'�5�)�W���	Ӊ��@%��Q*��'���u�u�u�u�>�3�Ϸ�Yђ��VD��N����� �0�>�0�w�;��������G��N��Oʦ�2�4�u�&�u�/���YӇ��A��C�����:�u���>�)�W���Y�����Y�����!� �w�_�w�)�����Ƨ�V��QN��6����!��9�w�}�W�������@F��E��N���4�!�<� �2�6����ӕ��\��R/�����9�o�&�2�6�}�������9F��C�����u�0�%�:�w�.�������F�T�����9�<�u�!�"��}�������F��\��U���&��0���$�W���Y�ƿ�T����W���0�n�_�u�#�/����Y����U��B����;�n�u�4�#�4��������R��CN��U���:�3�1�'�4�}�W�������@F�UךU���'�7�!�u�6�����Ӊ��@��R�����9�o�&�2�6�}����[���R��^��ʸ�-�3�;� �w�;��������TF�T�����9�<�u�m�l�W����s���F��P�����9�u�;� �$�)�W�������R��Y�����<�4�:�<�;�1�����Ƹ�VF��=N��Xʱ�4�'�8�u�u�8����Ӓ��@��^	�����:�4�:�1�:�/��������G��X���ߊu�x�3�9�2�.�����Ɖ��������:�0�:�u�?�.�W�������R��E��U���0�!�,�u�z�}�Ϫ�ӵ��C
��[��U���4�;�u��>�}��������V��qI�����4�9�!�u�?�}�W��Y����A��fN�����y�4�1�?�$�}����
Ӓ��
��S��U���!�0�6�0�1�>����Y���F�_�����{�u��2�$�8�6�������	l�G������8�9��<�W�W������F�������0�2�}�4�'�8��������F�N�����:�1�0�u�j�.��������F�N�����0�0�u�h�$�2����s���F��X�����2�i�u��2���ԜY�Ʃ�WF��d�����%�:�0�&��:����8����C��dךU����<�u�:�2�>����Y����[F��R�����!�"�r�0�8�}�GϪ�Y����A��T��\���;�u�u�x�w�<�W�������A��D��U���>�0�u�'�4�}�ϩ�����r%��RI��U���}�&�0�=�1�t�}�������@%��Y��O���%�:�0�&��0�������Q��Yd��Uʼ�u�<�<�2�2�:�_���	����XO��_�����u�u�3�&�8�;�������F��R ךU���u�u��0��(����E����G��DS�E���_�u�u�u�w�
�$������Z������k�e�|�_�w�}�W���.����U�N��H��r�_�u�u�w�1����:����V4��
I�U���;�u�u�u�w�4�W�������]��
�����:�>�d�!�2�W�W���Y���@%��Q-�����u�h�}�!�2�.�I��P���F�N�����=�3�u�h�$�8����Q����~��\�����:�e�u�u�g�f�W���Y����_��N��U���u�&�:�3�8�3����Dӕ��V ��B �����d�_�u�u�w�}�������F�R ����_�u�u�;�w�;�}����Ƽ�\��DN�����&�:�;�0�l�W�W�������g	��D�Uʥ�:�0�&��:�1�4������Q��Yd��Uʼ�u�<�<�2�2�:�_���	����X(�������u�u�&��2��������@��[�����6�:�}��2�������ƹF������;��0�&�4�}�Jϭ�����G]ǻN��U���:�3�0�i�w�����+����F�N��6�����,�i�w�.�������F��SN��N���0�1�%�:�2�.�#���
����\ ��CUװUʦ��0��1�w�`��������A*��d�����4�<�2�:�1�}�Jϭ�5����]��R����_�u�x�u�?�.����Y����@F��S�����u�'�!�u�9�?�����Ʃ�P��QN��ʘ��y�"�<�?�W�W��	������_N��ʺ�0�6�6�0�1�/����Y����U��R ��Uʚ�!� ��&�]�}����
�Ο�^��t���ߊu�0�<�_�w�}�Ϭ�
����V��=�����9��|�!�2�W�W���Y����zF��^��ʾ� ��6�x�w�2����Y�����X�����4��9��w�`��������p	��D"��]���4�1�&��2�
�W���Y����@��R��1���_�u�u�u�9�}����s���F��������2�r�r�#�8�}���Y���@��R�����9�i�u��2�����B���F��Y
���ߊu�u�;�u�1�W�W���Y����V��x�� ���&�_�u�&��8�3���Y����@%��Q*�����n�u�&��2�
�6��� ���@��R��4���,�6�n�_�9�}�#��