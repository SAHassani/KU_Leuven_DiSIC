-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����1�{�=�_�z�����CӬ��VF��Y�����u�'�2�;�;������Ɯ�z��Z������!�o�g�w�-����I��ƴl�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�u�4�}�G��:����Z�� �����9��&�'�:�3�ϝ�����G��=C�4����2�!�u�2�8����T�Ƃ�G��V����� �0�!�u�9�8����0����^��X חX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�Z�������V\�:��ʳ�9�u�;�!�9�4��������x��EN�>���<�%�0��6�}����;����R��V�����&�x�u�u�w�}�W�������V��[��ʡ�0�6�;�0�#�2�ϼ�������*��ʘ�8�'�u�;�w�5�W���4���F�N��U���0�:�'�0�w�3����?����9K��C��U���u�u�u��:�1�W���Ӷ��GF��v#��ʺ�0�:�u�=�w�2��������G��U�����-�7�:�>���}��Y���F�N��U�������w�5�����Ƹ�\F��S�����!�%�'�&�w�3�W���Ӗ��GF��SN��ʢ�<�0�x�u�w�}�W���YӖ��GH��Y��ʺ�=�'���w�2�������w6��e/�����u�9�:�&�"�}�Ͽ�N�Ʈ�GF��CחX���u�u�u�u�w�(�[ϼ�Y����A	��D��U���=�4�&�4�;�*���KӃ��^��DN����� �4�<�;�]�p�Z���Y���F�:��U���<�;�0�0�2�)����Y����[��v#�����{��u�4�w�/��������]��S��X���u�u�u�u�w�;�ψ�����F��p/��U���u�:�u�<�#�%�W���
����G��C��U���8�;�u�:�]�p�W���Y���F�������0�!���/�l����=�ơ�W�C��U���u�u�u���l�$����ƭ� P��^�����g�1�0�y�f�}�ϭ�����W����ʇ��_�x�u�w�}�W���Y���� P��gN��U���g�7�!�7�w�l�W���	����-��D����� �9�%�'�w��Y��s���F�N��Uʂ�<�<�2�!�8��W���	����Z��CN��ʦ�8�u�<�0�>�}��������3�������,�<�0�x�w�}�W���Y����\F��R��ʡ�0�&�/�u�1�)�Ϻ��Ʈ�@HǶd�U���u�u�u�u��8�8����ƞ�T��R��ʡ�0���u�$�8����Ӏ����C�����{�x�u�u�w�}�W���-����Z��^ �����,�7�!�0�9�.��������@F��SN����� �u�&�g�4�>���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����'�'�u����}���
�ƙ�z5�������0�!�{�9�l�1���� ӳ��~'��xUךU���u�����+����������d�����'�u�0�0�w�2��ԜY����Z����*���<�
�d�a�6�1�}���
�ƥ�V��B�����!�{�9�n�w�(�ϩ��Ȝ�T(��C������%�4�9�]�}��������X��G@���ߠ0�!�!�u�%�>�3�������CF��=N�����<�}�u�u�<�<����*����\��YN�����'�'�;�0�f�)�W���C����l�G��]���u��8�9��6�W���Cӏ��@��[���ߠu�u�&�'�#�����
����]F��D�����u�:�;�:�g�f�W���
����z��[��U���;��:�0�9�8��������r��^��X��1�"�!�u�~�W�W���=����]/�N��Oʼ�u�<�;�1�o�/����Q����R'��d��U���u�:�;�:�g�f�Z���H����F�D*�����u�u�u�o�>�}�����ލ�A��CF�����'��/�u�w�}�������K�d_�D�ߊu�u��4��9����Y�ƥ�F��D�����u�:�;�:�g�f�W���
����|��N��U��� �u�<�;�3�e����&�Χ�R��E�����u�u�:�;�8�m�L��Y����l�N����� ��u�u�m�2�ύ�����'��V��]���!��,�<�2�p�FϺ�����O�C�&��d�_�;�u�%�>�3�������C]ǑV�����!�'�u��w�;�1�������A��S���ߊu�:�%�;�9�}�6���O����F�P�����}�u�u�u���2���Y���F�N��U���0�0�u�u�w�`�G�ԜY���v(��t-��0���u�u�u�u�m�?�������\�q/��0�ߊu�u�u����$���;���F�N�����;�u�u�o�w��$��Y���#��r-��"����u�u�u�w�}�������F��(��&��u�u�u���}�W���Y���F�T�����0�!�'�u�j��G��I����V��^�E��u�u�u����>���Y���F�T�����2�u�u�u�j��8���B���F��~#��:�����
���}�W������F�S��4���n�u�u�u���:���Y���F�N��U���<�2�u�u�w�`�U���<��ƹF�=��4���u�u�u�u�w�}�W�������P��N�U���e�e�e�e�g�m�G��I����F�G��U�ߊu�u�u����W����ƿ�W9��X	��N���u�u��u�w�(�W���&����P9��T��]��1�"�!�u�~�W�W���Y����	F��CN�����2�6�#�6�8�u�W������]ǻN��U������u�w�(�W���&����P9��T��]���:�;�:�e�l�}�W���*����a4���U���
�9�2�6�]�}�W���=����Z��C
�����
�0�!�'�a�}�������9F�N��<���u�;�&�1�;�:��������F��@ ��U���_�u�u�u���%���ƿ�W9��P�����:�}�u�:�9�2�G��Y���4��{%��U���&�1� �:�>�f�W���YӴ��}F��^ �����9�2�6�_�w�}�W���:����Z��C
�����6�_�u�u�w��W���ӕ��l��P�����u�u��o�>�}��������E��X��U���;�:�e�n�w�}�Wω�8����	F����*���<�
�0�!�%�e��������l�N��"����o�<�u�#��������F�`<��U���;�&�1� �8�4�^�ԜY����P	��X ���ߠu�6�8�:�2�)�%���H˵��9F�	�����u�_�u�u�w��%���Y���F�N��Oʼ�!�2�'�u�w�g�W��Y���/��cN��U���u�u�u�u�w�}��������F��6��E��e�e�e�e�g�m�G��Y���/��c1��9���u�u�u�u�w�}�������F��L��;���_�u�u�u���8���*����p.��|N����;�u�u�u�m�}�6���B���F��~#��:���u�u�u�u�w�}�W������F�S��&���w�_�u�u�w��6���Y���F�N��Oʷ�!�#�6�:�w�g�W���I����V��^�E��w�n�u�u�'�/�W�ԜY���w)���U���
�:�<�
�2�)���Y����G	�UךU���u��u�u�"�}��������E��X��U���;�:�e�n�]�}�W���0����]F��S1�����#�6�:�}�f�9� ���Y����F�N��%��<�u�!�
�8�4�(��������Y��E��u�u�u����W���ӕ��l
��^�����'�m�1�"�#�}�^�ԜY���a"��|N����!�
�9�2�4�W�W���Y����\��YN�����:�<�n�u�w�}�%���<����]F��S1�����n�u�u�u���MϷ�Y����F
��^�U���u��u�u�9�.��������V��EF����!�u�|�_�w�}�W���=�����D�����6�#�6�:��}�������9F�N��'���u�u�;�&�3�(����B���F��e+��Oʼ�u�!�
�9�0�>�L�������\��Y��N�ߊu�u�x��2��6�������R������7�!�4�1�2�.�}���Y����R
��z�����'�o�&�1�;�:��������F��@ ��U���h�}�!�0�$�`�W��P���F��P ��U���8�1�1�'�m�.��������V��EF����!�u�|�h��)����D���O��=N��U����0�����W���Y����C��R ��W���0�"�1�w� �4�ϻ�����l�N�U���=��u�:�#�2�ϱ�ӄ��VF��*�����:�0�7�!�8�}�>��Y���F�� ��ʡ�u�9�6�u�?�}��������
K��CN�����u�=�!�&�6�8�ω�s���K��XN�����<�1�%�;�2�)� ����ƪ�AF��T��$ʦ�8�9�{�u�w�>�����Ƨ�V1��C��1����&�u�o�>�)����C����9F������!�>�0�<�#��'�������\��Y�����h�d�_�u�w�2����Ӎ��d��_N��U���u�u�u�u�9�8����DӍ��d��_!����� �~���3�5��������@]ǑN��X����&�8�9�$�<���Y����D��N�����4�%�0�<�w�<��������Q��Dd��U���u�;��z��<�������\��~>��:�ߊu�u�:�&�6�)��������[F��^ �����o�u�m�_�w�}��������z��Z��"���=�o�<�!�0�/�M���=����Z��\�U���6�;�!�;�w���������A5��G��Oʼ�!�2�'�o�w��$�������G��`�����_�u�u�!�'�}��������E9��^�����}��!��.�4���Hӂ��]��G��ʦ�1�9�2�6�!�>����0����C
��^
��X���:�;�:�e�l�}�Wϭ�����@"��V'�����u�u�4�4�9�,����B���F������<�&�0��:�1�W����Ƽ�AF��Z��[���u�!�%�u�2��6���ӏ��R��NF�����'��/�x�w�2����I�ƣ���h�����0�!�'�>�2�4����=����F��z�����&�0��8�;�p�W������]ǻN�����9�&�0���$�Mϓ�����J9��=N��U���;�9�&�0��}�W���&����P9��T��]����1�=�;�6�<����4����q��g�����0�>�4�4�%�����Y�ƨ�D��^����u�<�;�9�$�8�3���Y����_	��T1�����}���1�?�3�����̧�V��u��%���4�%�0�>�6�<�������F��@ ��U���_�u�u�<�9�1��������B'��q��U���!�
�:�<��8��������^��`�����4�4�'��-�}�W�������V�=d��U���u��8�0�>�.��������Q����U���%�0�u��%�)�W���
Ӈ����SN��U���4�_�u�u�.�8�:�������l��DN�����>�4�4�'��'�Z�������V�X�����:�<�
�0�#�/��������]6��^�� ����8�0�<�$�8�$�������W	��C��\�ߊu�u�<�;�;�.����	����	F��Z*��4���!�_�u�u�>�3�ϭ�����\��C
�����
�0�!�'�<�8����6����Z��B��8���0�<�&�0��0����=����A��M��U���:�;�:�e�l�}�Wϭ�����@+��s!��Oʦ�1�9�2�6�!�>����.����G��g�����&�>�0���)�'���������C�����0�x�d�1� �)�W���s���K�c��"���'�4�{�u�w�.����Y����d��NN����9�2�6�#�4�2�_�������G��E=�����>�4�4�'��'�W���Y����G	�UװUʷ�2�;�_�u�w�8� �������R0��^
���ߊu�u�:�u�w�3��������Z��N�����u�u�0�0�6�8�W���Y���p��C������4�'�,�1�/��������JHǻN��U����6�u��$�0����
����~��R,������8�9�u�6�<����
Ӈ����^�����{�u�u�u�z�}�ϰ��Ƹ���[
��ʴ�'�,�!�4�w�2����
Ӄ��[F��V�����<�u�:�u�w�}�Z���4����q��g�����0�0�0�0�#�}�Ϫ�ӕ��^1��E�U���u�&�0���$����.����@6��d�����<�d�u�u�w�2��������V$��D>��&���9��|�i�w�2����Y����\9��S������!���;�9����B�����	�����0��;�0�%�0��������A��=N��U����;�0�!�#�8����Y����D��RN�����&�&�_�u�w��������F��S1�����#�6�:�}� �4��������l�N������1�u�h�$�9��������G	��D<�����'�&�|�_�w�}�0�������`
��=N��U���u�u�;�>�6�<�������F��@ ��U���0�0�4�0�w�}�W��Y����C��QN�����!�u�<�&�6�8��������G	���ʺ�u��4�1�f�?�ϱ�Y����9F�N��1������#�>�}�Jϭ�����Z��R��¦�4�4�;�}�~�}�W���&����P9��T��]���!���<�~�W�W���YӶ��X+��s��O���u�u�3�'�=�4�W�������G��E=�����x�d�1�"�#�}�W�������9F�N��U����:�%�u�1�6�����Ʈ�G��E�����;�1�!�u� �
��������G��DN�����;���4�3�6��������R��B�����:�u��_�w�}�W���4����C'����]����1�=�;�6�4����P�Φ�O�_�����:�}���3�5��������@O��N�U���!����!�4�_���.����N��G��U���:�;�:�>�2�4�������F��R9������'�!��$�f�W���Y����~��^/��U¼�}�>�0�<�#��3���;���L��_��X��1�"�!�u�<�8����6����R$��N�����h�&�4�4�9�,����Pۍ��d��_D��^ʾ�0�<�!���)�5���T����\��XN�����!��|�_�w�}�W���Y����A��>������!�n�u�w�8�Ϲ�����VF��Y'�����9�n�_�u�w�8�Dٕ�;����W��N��X���0�0�!�!�2�.����Ӓ����X�����;�<�2�:�w�2�W��� Ӗ��R
��[N�����&�4�0�'�&�4���Y����UF��V�����/�u�u�u�2�8����Y���K�q�����!�0�&�0���Ͽ�ӕ��^"��v��U���u�&�0��w�a�W�������JN��N�������,�e�l�}�W���
����z6�
N�����%�'�}�|�q�.����	����O��=N��U�����c���}�W���;�П�cl�N��Uʲ�;�'�6�8�'�W�W���Y���w)��r)��U���u�u�u�u�j�}�[���Y���F��y1��6����u�u�u�w�}�Iϸ�����F�N��Uʐ�
��
���}�W���Y���U��RBךU���u�u�u�x��/�W���Y����v%��R �����<�u�=�u���W���
ӏ��A��^��U��� �0�!�0�'�/��ԜY���F�C�����4�u�4�4�]�}�W���Y�Ɖ�l#��h9��!���u�u�u�h�w�<���Y���F�'��!���u�u�u�u�w�}�W���!����V��^�E��e�e�y�u�w�}�W���0����u/��N��U���u�u�k�w���[���Y���F��~#��:�����
���}�I���5����9F�N��U����
���w�}�W���Y���D��q+�����u�u�u�u���W���Y���F�N��U���e�e�e�e�g�m�G��I��ƹF�N�����8�%�_�u�w�}�W���TӲ��#��X�����6�<�;��3�}�2���Y����\��D�����u�u�u�u���%���Y����C��=N��U���u�u����}�W�������9F�N��U������u�w�c����U���F�N��X��� �%�!�'�0�.����
����A	��B�����{��!� �2�s�W���Y���5��S�R��_�u�u�u�w�}�Z�������c	��=N��U���u�u���w�`�W���	����XJǻN��U���u��u�u�j�}�:�������9F�N��U������h�w���������F�N��Uʑ�u�u�u�k�$�8�3��Y���F�*��U���h�u��8��q�}���Y���F�9��;���'�!�u�:�#�����P���F�N��X���=�u�'�!�w�2�Ϸ�Y����_��V�����!�8�{�u�w�}�W���T�ƛ���B��U���&�%�:�!�$�3����������C�����u�u�u�u���W��Y���9l�N��U���x�u�0�1��/�}���Y���F��t"��U���8�9��<�W�W���Y���a"��N��K��r�u�x��6�}�����Ƙ�VF��V
�����<�u�;�7�2�}�����Ƹ�^�N��U���u����w�c�P���Y����F��CN�����0�&�0�4�;�9�}���Y���F��v*��U��&�0���3�q�W���Y���"��N��H����8��_�w�}�W���Y����F�	N������n�u�u�2�9��������t��%�����1�n�_�u�w�8�Fו�;����W��N������!��,�>�8�J������R��N��U���u�&�<�;�#�8����=������������,�!�u�w�)�(�������P��d��U���&�0��u�k�}�:�������O��N��Uʦ�0���i�w�����8���]ǑN��Uʇ��d���/�g�%���H˵��9F�N��U���0�<�u�4��}�W���Y����|9��pN��U���u�u�u�u�i�l�}���Y���F��~:��U���u�u�u�u�w�`�W���I����V��^�E��w�_�u�u�w�}�W���-����vF�N��U���h�u���u�W�W���Y���`/��t!��<�������j�}�6���U���F�N��<�����u�u�w�}�W���G�ğ�u#�=N��U���u�u���w�}�W���Y���F�6��E��e�e�e�e�g�m�G���Y���F�C�����u���m��}��������R��r-�����9�7�0�_�w�}�W�������R�N��U���u�x�u� �'�)����
������T�����u�0�0�{��)����W���F�N��&���u�u�u�k�p�z�}���Y���F�N������'�_�u�w�}�W���+����[�d�����>�_�u�u�w�}�W���Y���F��R��4���_�u�u�u�w�}�%���+���@+��`�����u�u�u�u�w��W���Y����~��~BךU���u�u�u��w�}�J���4����cJǑN��U���u�x�u���u����Y����#��U��[���u�u�u�u�z�}��������C	�������9�1�4�9�#�8����W���F�N��Xʂ�u�&� �0�w�2��������Z��RN�����u�'�!�&�]�}�W���Y�ƛ�v(�S�R��_�u�u�u�w�}�Z�������\��N��U���u����w�c�$�������l�N��U�����u�u�i�z�P���TӴ��WF��V��[ʁ�0�'�4�u�8�)��������WF��[N��ʡ�8�{�u�u�w�}�Wό�>���X�I�X��� �%�!�'�0�.��������V�N��U���u����w�c����+����AJǻN��U���u��u�u�j�}�:���6���F�N��1���u�u�k�&�2��'��Y����]��R ������;�m�7�%�0���s���f��T�����4�_�u�u�8�}�W�������r��^�������!��%�<����T����\��XN����'�!�_�u�w�}�Zό�����]F��RN��U���0�u�;�u��}�����Ɓ�^"��V!��U���2�:�%�u�1�6�����Ʈ�G�N��Uʦ�4�4� ���$��������W����\���d�1�"�!�w�
� ����Υ�O���"���=�;�4�<�.�(�^��Y����w)��\9�������'�!��.�_���P�����Y�����<�!���%�)�5�����ƹF������!�$�'��6�u� �������M��`�����;�4�4� �w�l�����Ƨ�V1��C��\���u�u�u�u�w�`����=�Χ�V1��C��1����&�}�~�~�p�FϺ�����X1��^
��:���!��&�<�l�}�Wϻ�Ӂ��V��RN������8�4�4�]�}�Z���
�����������u�;�:�4�$�:��������9F��R �����!�'�o�u�w�;�Ϸ��Ƨ�R��E�����u�u�:�;�8�m��������F�D*������<�u�h�$�:����=����F��v�����>�$�4�%�2�4�������F��S�������8�9� �9�ŷ�RӍ��G��S��\�ߊu�u��!��)�_���E�ƿ�T�������!�$�'��6�u�>�������Z����U���!��1�=�z�l�����Ƨ�B5��G������|�n�u�2�9��������t��V�� ���,�_�;�u��f