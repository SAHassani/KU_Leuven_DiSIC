-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B"��V#�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������4ǶN����g�u�0�0�5�/�E��s��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�}�|�e�l�W��� ����GF��C�����;�!� �0�#�}��������]l�/��U���=�&��&�%�8�}��7����]��~ �����;�&��!�%�<�W�������Z	��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�'�������g�������;�u�8�9�:�3�Ͽ�����d��_N�����%�!�u�u�2�-�W���T����WFǶN�����!�'�2�&�2�s�W���Y����Z��YN�����u�;�,�6�9�/��������TF��C��ʡ�0�x�u�u��q��������F��CN��[����!��1�?�4�W�������W����U���u�0�&�!�]�p�W϶�����Z ��R�����x�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s���Q��NN����u� �0�<�2�s��������W����N��� �0�<�0�y�(����&����R
��=d�U���!�0�<�u�%�3����&������V��-���;��'��5�W�����ƙ�z5��d��ʀ���{�6�:�2����W����9K�D�����&�!�4�&�6�8��Զs����G��F*�����:�,�<�u�]�8����Q����w��`�����u�u�;�<�#�:���s����l�d�����>�-�u�o�>�}��������9F��D*�����u�u�u�u�9�.��������V��EF�����<�!�x�u�8�3���B����@1��C��U���u�u�;�&�3�1����s�ƿ�r��R��U���o�<�u�!��2��������W��X����n�u�&��#�����Y����F��C
�����
�0�!�'�<�<��������W	��C��\���_�;�u�$�6�<���� ��ƓR��^�����u��u�3����������ZǑN�����0�!���d��W���	����l�N�����o�<�u�!��2����D����l�N����<�u�!�
�8�4�W��^����F�N��U���;�&�1�9�0�>�M���I��ƹF���U���&�1�9�2�4�+����Q�ƨ�D��^����u�u�u�u�"�}��������9F�N��F���u� �u�!��2����s�Ʃ�WF��Z�����_�u�x�=�8�������ƹK��_��*���0�1�_�u�>�3�ϭ�8����@��[��U���
�:�<�
�2�)�������\F��N��U���u�u�o�u�8�5���^���9F��^	��ʦ��!��!�8�?�Mϭ�����Z��R��¾�4�4�<�!�z�}�������	[�X����r�r�n�u�$�:����
����|��T��Oʦ�1�9�2�6�!�>����=����Z��_�����:�e�u�h��)����G���l��R	�����&��1�0�$�(���Y����F�D�����&�_�u��9���ԜY����zF��^��ʾ�4�4�<�!�z�}������ƹF��������g�_�w�}�Z�������P
��d�����>�-�u�u�z�+����ӂ��@"��V'��<�ߊu�u�x�=�8��W���
����G��=N��U���=�:�
�u�w�.����
����_l�N����>�4�$�&��)�8�������l�N����>�4�$�d�8�8�}���Y���� T��N��9���u�u�u�'�/�W���Y���F�N����u�4�%�0�;��[���Y���F��N�����2�6�o�u�g�W�W���Y�ƨ�F������;��y�u�w�}�Z����ƿ�W9��P��O���e�_�u�u�w�}����Gӕ��A��r �U���u�u�x�u�9�}��������	[�IךU���u�u�u�u�i�.�6�������_
�N��X���;�u�!�
�8�4�(��������Y��E�ߊu�u�u�u�w�}�Iϭ�=����F��Z��\���x�u� �u�#�����s���F�F]�H���%�;�n�u�w�}�W���Y���\��D�����6�u�0�1�0�3����Y����a*��=d��3���9�3�_�u�%�>��������p
��OGךU���<�_�u�u�1�/����&����5��G�����|�!�0�_�w�}�W�������G*��R�����!��!�:�5�W�W����ƥ�l�R �����0�&��;�;�;�}���
����R)��R�����!��!�6�l�W����-���